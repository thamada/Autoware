-- ==============================================================
-- Time-stamp: <2017-01-04 22:08:27 hamada>
-- Copyright (C) 2017 Tsuyoshi Hamada. All Rights Reserved.
--
-- Autoware for FPGAs project.
-- 
-- --------------------------------------------------------------
-- RTL design for my OpenCL-enebled custom GPU
-- ==============================================================

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gpu is
generic (
    C_M_AXI_GMEM_ADDR_WIDTH : INTEGER := 32;
    C_M_AXI_GMEM_ID_WIDTH : INTEGER := 1;
    C_M_AXI_GMEM_AWUSER_WIDTH : INTEGER := 1;
    C_M_AXI_GMEM_DATA_WIDTH : INTEGER := 32;
    C_M_AXI_GMEM_WUSER_WIDTH : INTEGER := 1;
    C_M_AXI_GMEM_ARUSER_WIDTH : INTEGER := 1;
    C_M_AXI_GMEM_RUSER_WIDTH : INTEGER := 1;
    C_M_AXI_GMEM_BUSER_WIDTH : INTEGER := 1;
    C_S_AXI_CONTROL_ADDR_WIDTH : INTEGER := 7;
    C_S_AXI_CONTROL_DATA_WIDTH : INTEGER := 32;
    C_M_AXI_GMEM_CACHE_VALUE : INTEGER := 3;
    C_M_AXI_GMEM_USER_VALUE : INTEGER := 0;
    C_M_AXI_GMEM_TARGET_ADDR : INTEGER := 0;
    C_M_AXI_GMEM_PROT_VALUE : INTEGER := 0 );
port (
    ap_clk : IN STD_LOGIC;
    ap_rst_n : IN STD_LOGIC;
    m_axi_gmem_AWVALID : OUT STD_LOGIC;
    m_axi_gmem_AWREADY : IN STD_LOGIC;
    m_axi_gmem_AWADDR : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_ADDR_WIDTH-1 downto 0);
    m_axi_gmem_AWID : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_ID_WIDTH-1 downto 0);
    m_axi_gmem_AWLEN : OUT STD_LOGIC_VECTOR (7 downto 0);
    m_axi_gmem_AWSIZE : OUT STD_LOGIC_VECTOR (2 downto 0);
    m_axi_gmem_AWBURST : OUT STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem_AWLOCK : OUT STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem_AWCACHE : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem_AWPROT : OUT STD_LOGIC_VECTOR (2 downto 0);
    m_axi_gmem_AWQOS : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem_AWREGION : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem_AWUSER : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_AWUSER_WIDTH-1 downto 0);
    m_axi_gmem_WVALID : OUT STD_LOGIC;
    m_axi_gmem_WREADY : IN STD_LOGIC;
    m_axi_gmem_WDATA : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_DATA_WIDTH-1 downto 0);
    m_axi_gmem_WSTRB : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_DATA_WIDTH/8-1 downto 0);
    m_axi_gmem_WLAST : OUT STD_LOGIC;
    m_axi_gmem_WID : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_ID_WIDTH-1 downto 0);
    m_axi_gmem_WUSER : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_WUSER_WIDTH-1 downto 0);
    m_axi_gmem_ARVALID : OUT STD_LOGIC;
    m_axi_gmem_ARREADY : IN STD_LOGIC;
    m_axi_gmem_ARADDR : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_ADDR_WIDTH-1 downto 0);
    m_axi_gmem_ARID : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_ID_WIDTH-1 downto 0);
    m_axi_gmem_ARLEN : OUT STD_LOGIC_VECTOR (7 downto 0);
    m_axi_gmem_ARSIZE : OUT STD_LOGIC_VECTOR (2 downto 0);
    m_axi_gmem_ARBURST : OUT STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem_ARLOCK : OUT STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem_ARCACHE : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem_ARPROT : OUT STD_LOGIC_VECTOR (2 downto 0);
    m_axi_gmem_ARQOS : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem_ARREGION : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem_ARUSER : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_ARUSER_WIDTH-1 downto 0);
    m_axi_gmem_RVALID : IN STD_LOGIC;
    m_axi_gmem_RREADY : OUT STD_LOGIC;
    m_axi_gmem_RDATA : IN STD_LOGIC_VECTOR (C_M_AXI_GMEM_DATA_WIDTH-1 downto 0);
    m_axi_gmem_RLAST : IN STD_LOGIC;
    m_axi_gmem_RID : IN STD_LOGIC_VECTOR (C_M_AXI_GMEM_ID_WIDTH-1 downto 0);
    m_axi_gmem_RUSER : IN STD_LOGIC_VECTOR (C_M_AXI_GMEM_RUSER_WIDTH-1 downto 0);
    m_axi_gmem_RRESP : IN STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem_BVALID : IN STD_LOGIC;
    m_axi_gmem_BREADY : OUT STD_LOGIC;
    m_axi_gmem_BRESP : IN STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem_BID : IN STD_LOGIC_VECTOR (C_M_AXI_GMEM_ID_WIDTH-1 downto 0);
    m_axi_gmem_BUSER : IN STD_LOGIC_VECTOR (C_M_AXI_GMEM_BUSER_WIDTH-1 downto 0);
    s_axi_control_AWVALID : IN STD_LOGIC;
    s_axi_control_AWREADY : OUT STD_LOGIC;
    s_axi_control_AWADDR : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_ADDR_WIDTH-1 downto 0);
    s_axi_control_WVALID : IN STD_LOGIC;
    s_axi_control_WREADY : OUT STD_LOGIC;
    s_axi_control_WDATA : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_DATA_WIDTH-1 downto 0);
    s_axi_control_WSTRB : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_DATA_WIDTH/8-1 downto 0);
    s_axi_control_ARVALID : IN STD_LOGIC;
    s_axi_control_ARREADY : OUT STD_LOGIC;
    s_axi_control_ARADDR : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_ADDR_WIDTH-1 downto 0);
    s_axi_control_RVALID : OUT STD_LOGIC;
    s_axi_control_RREADY : IN STD_LOGIC;
    s_axi_control_RDATA : OUT STD_LOGIC_VECTOR (C_S_AXI_CONTROL_DATA_WIDTH-1 downto 0);
    s_axi_control_RRESP : OUT STD_LOGIC_VECTOR (1 downto 0);
    s_axi_control_BVALID : OUT STD_LOGIC;
    s_axi_control_BREADY : IN STD_LOGIC;
    s_axi_control_BRESP : OUT STD_LOGIC_VECTOR (1 downto 0);
    interrupt : OUT STD_LOGIC );
end;


architecture behav of gpu is 
    attribute CORE_GENERATION_INFO : STRING;
    attribute CORE_GENERATION_INFO of behav : architecture is
    "gpu,hls_ip_2016_4,{HLS_INPUT_TYPE=c,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcku025-ffva1156-1-c,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=8.750000,HLS_SYN_LAT=551,HLS_SYN_TPT=none,HLS_SYN_MEM=2,HLS_SYN_DSP=2,HLS_SYN_FF=2015,HLS_SYN_LUT=2034}";
    constant ap_const_logic_1 : STD_LOGIC := '1';
    constant ap_const_logic_0 : STD_LOGIC := '0';
    constant ap_ST_fsm_state1 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
    constant ap_ST_fsm_pp0_stage0 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
    constant ap_ST_fsm_state139 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100";
    constant ap_ST_fsm_pp1_stage0 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000";
    constant ap_ST_fsm_state277 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000";
    constant ap_ST_fsm_state278 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000";
    constant ap_ST_fsm_state279 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000";
    constant ap_ST_fsm_state280 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000";
    constant ap_ST_fsm_state281 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000";
    constant ap_ST_fsm_state282 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000";
    constant ap_ST_fsm_state283 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000";
    constant ap_ST_fsm_state284 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000";
    constant ap_ST_fsm_state285 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000";
    constant ap_ST_fsm_state286 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000";
    constant ap_ST_fsm_state287 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000";
    constant ap_ST_fsm_state288 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000";
    constant ap_ST_fsm_state289 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000";
    constant ap_ST_fsm_state290 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000";
    constant ap_ST_fsm_state291 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000";
    constant ap_ST_fsm_state292 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000";
    constant ap_ST_fsm_state293 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000";
    constant ap_ST_fsm_state294 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000";
    constant ap_ST_fsm_state295 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000";
    constant ap_ST_fsm_state296 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000";
    constant ap_ST_fsm_state297 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000";
    constant ap_ST_fsm_state298 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000";
    constant ap_ST_fsm_state299 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000";
    constant ap_ST_fsm_state300 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000";
    constant ap_ST_fsm_state301 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000";
    constant ap_ST_fsm_state302 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000";
    constant ap_ST_fsm_state303 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000";
    constant ap_ST_fsm_state304 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000";
    constant ap_ST_fsm_state305 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
    constant ap_ST_fsm_state306 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000";
    constant ap_ST_fsm_state307 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000";
    constant ap_ST_fsm_state308 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000";
    constant ap_ST_fsm_state309 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
    constant ap_ST_fsm_state310 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000";
    constant ap_ST_fsm_state311 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000";
    constant ap_ST_fsm_state312 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000";
    constant ap_ST_fsm_state313 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000";
    constant ap_ST_fsm_state314 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000";
    constant ap_ST_fsm_state315 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state316 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state317 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state318 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state319 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state320 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state321 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state322 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state323 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state324 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state325 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state326 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state327 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state328 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state329 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state330 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state331 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state332 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state333 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state334 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state335 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state336 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state337 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state338 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state339 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state340 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state341 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state342 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state343 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state344 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state345 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state346 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state347 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state348 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state349 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state350 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state351 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state352 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state353 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state354 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state355 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state356 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state357 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state358 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state359 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state360 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state361 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state362 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state363 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state364 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state365 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state366 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state367 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state368 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state369 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state370 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state371 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state372 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state373 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state374 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state375 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state376 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state377 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state378 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state379 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state380 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state381 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state382 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state383 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state384 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state385 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state386 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state387 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state388 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state389 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state390 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state391 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state392 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state393 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state394 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state395 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state396 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state397 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state398 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state399 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state400 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state401 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state402 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state403 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state404 : STD_LOGIC_VECTOR (143 downto 0) := "000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state405 : STD_LOGIC_VECTOR (143 downto 0) := "000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state406 : STD_LOGIC_VECTOR (143 downto 0) := "000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state407 : STD_LOGIC_VECTOR (143 downto 0) := "000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state408 : STD_LOGIC_VECTOR (143 downto 0) := "000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state409 : STD_LOGIC_VECTOR (143 downto 0) := "000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state410 : STD_LOGIC_VECTOR (143 downto 0) := "000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state411 : STD_LOGIC_VECTOR (143 downto 0) := "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state412 : STD_LOGIC_VECTOR (143 downto 0) := "000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state413 : STD_LOGIC_VECTOR (143 downto 0) := "000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state414 : STD_LOGIC_VECTOR (143 downto 0) := "001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state415 : STD_LOGIC_VECTOR (143 downto 0) := "010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state416 : STD_LOGIC_VECTOR (143 downto 0) := "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_const_lv32_0 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000000";
    constant ap_const_lv1_1 : STD_LOGIC_VECTOR (0 downto 0) := "1";
    constant ap_const_lv32_1 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000001";
    constant ap_const_lv1_0 : STD_LOGIC_VECTOR (0 downto 0) := "0";
    constant ap_const_lv32_3 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000011";
    constant ap_const_lv32_5 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000101";
    constant ap_const_lv32_C : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001100";
    constant ap_const_lv32_8F : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000010001111";
    constant C_S_AXI_DATA_WIDTH : INTEGER range 63 downto 0 := 20;
    constant C_M_AXI_DATA_WIDTH : INTEGER range 63 downto 0 := 20;
    constant ap_const_lv32_4 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000100";
    constant ap_const_lv32_6 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000110";
    constant ap_const_lv32_7 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000111";
    constant ap_const_lv32_B : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001011";
    constant ap_const_lv32_2 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000010";
    constant ap_const_lv5_0 : STD_LOGIC_VECTOR (4 downto 0) := "00000";
    constant ap_const_lv32_10 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000010000";
    constant ap_const_lv3_0 : STD_LOGIC_VECTOR (2 downto 0) := "000";
    constant ap_const_lv2_0 : STD_LOGIC_VECTOR (1 downto 0) := "00";
    constant ap_const_lv4_0 : STD_LOGIC_VECTOR (3 downto 0) := "0000";
    constant ap_const_lv4_F : STD_LOGIC_VECTOR (3 downto 0) := "1111";
    constant ap_const_lv32_8 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001000";
    constant ap_const_lv32_1F : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000011111";
    constant ap_const_lv5_10 : STD_LOGIC_VECTOR (4 downto 0) := "10000";
    constant ap_const_lv5_1 : STD_LOGIC_VECTOR (4 downto 0) := "00001";
    constant ap_const_boolean_1 : BOOLEAN := true;

    signal ap_rst_n_inv : STD_LOGIC;
    signal ap_start : STD_LOGIC;
    signal ap_done : STD_LOGIC;
    signal ap_idle : STD_LOGIC;
    signal ap_CS_fsm : STD_LOGIC_VECTOR (143 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
    attribute fsm_encoding : string;
    attribute fsm_encoding of ap_CS_fsm : signal is "none";
    signal ap_CS_fsm_state1 : STD_LOGIC_VECTOR (0 downto 0);
    attribute fsm_encoding of ap_CS_fsm_state1 : signal is "none";
    signal ap_ready : STD_LOGIC;
    signal group_id_x : STD_LOGIC_VECTOR (31 downto 0);
    signal group_id_y : STD_LOGIC_VECTOR (31 downto 0);
    signal group_id_z : STD_LOGIC_VECTOR (31 downto 0);
    signal global_offset_x : STD_LOGIC_VECTOR (31 downto 0);
    signal global_offset_y : STD_LOGIC_VECTOR (31 downto 0);
    signal global_offset_z : STD_LOGIC_VECTOR (31 downto 0);
    signal x : STD_LOGIC_VECTOR (31 downto 0);
    signal y : STD_LOGIC_VECTOR (31 downto 0);
    signal z : STD_LOGIC_VECTOR (31 downto 0);
    signal x0_address0 : STD_LOGIC_VECTOR (3 downto 0);
    signal x0_ce0 : STD_LOGIC;
    signal x0_we0 : STD_LOGIC;
    signal x0_d0 : STD_LOGIC_VECTOR (31 downto 0);
    signal x0_q0 : STD_LOGIC_VECTOR (31 downto 0);
    signal y0_address0 : STD_LOGIC_VECTOR (3 downto 0);
    signal y0_ce0 : STD_LOGIC;
    signal y0_we0 : STD_LOGIC;
    signal y0_d0 : STD_LOGIC_VECTOR (31 downto 0);
    signal y0_q0 : STD_LOGIC_VECTOR (31 downto 0);
    signal gmem_blk_n_AR : STD_LOGIC;
    signal ap_CS_fsm_pp0_stage0 : STD_LOGIC_VECTOR (0 downto 0);
    attribute fsm_encoding of ap_CS_fsm_pp0_stage0 : signal is "none";
    signal ap_enable_reg_pp0_iter1 : STD_LOGIC := '0';
    signal isIter0_reg_481 : STD_LOGIC_VECTOR (0 downto 0);
    signal gmem_blk_n_R : STD_LOGIC;
    signal ap_enable_reg_pp0_iter135 : STD_LOGIC := '0';
    signal exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter134_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_CS_fsm_pp1_stage0 : STD_LOGIC_VECTOR (0 downto 0);
    attribute fsm_encoding of ap_CS_fsm_pp1_stage0 : signal is "none";
    signal ap_enable_reg_pp1_iter1 : STD_LOGIC := '0';
    signal isIter_reg_494 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_enable_reg_pp1_iter135 : STD_LOGIC := '0';
    signal exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter134_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal gmem_blk_n_AW : STD_LOGIC;
    signal ap_CS_fsm_state278 : STD_LOGIC_VECTOR (0 downto 0);
    attribute fsm_encoding of ap_CS_fsm_state278 : signal is "none";
    signal gmem_blk_n_W : STD_LOGIC;
    signal ap_CS_fsm_state285 : STD_LOGIC_VECTOR (0 downto 0);
    attribute fsm_encoding of ap_CS_fsm_state285 : signal is "none";
    signal gmem_blk_n_B : STD_LOGIC;
    signal ap_CS_fsm_state416 : STD_LOGIC_VECTOR (0 downto 0);
    attribute fsm_encoding of ap_CS_fsm_state416 : signal is "none";
    signal gmem_AWVALID : STD_LOGIC;
    signal gmem_AWREADY : STD_LOGIC;
    signal gmem_WVALID : STD_LOGIC;
    signal gmem_WREADY : STD_LOGIC;
    signal gmem_WDATA : STD_LOGIC_VECTOR (31 downto 0);
    signal gmem_ARVALID : STD_LOGIC;
    signal gmem_ARREADY : STD_LOGIC;
    signal gmem_ARADDR : STD_LOGIC_VECTOR (31 downto 0);
    signal gmem_RVALID : STD_LOGIC;
    signal gmem_RREADY : STD_LOGIC;
    signal gmem_RDATA : STD_LOGIC_VECTOR (31 downto 0);
    signal gmem_RLAST : STD_LOGIC;
    signal gmem_RID : STD_LOGIC_VECTOR (0 downto 0);
    signal gmem_RUSER : STD_LOGIC_VECTOR (0 downto 0);
    signal gmem_RRESP : STD_LOGIC_VECTOR (1 downto 0);
    signal gmem_BVALID : STD_LOGIC;
    signal gmem_BREADY : STD_LOGIC;
    signal gmem_BRESP : STD_LOGIC_VECTOR (1 downto 0);
    signal gmem_BID : STD_LOGIC_VECTOR (0 downto 0);
    signal gmem_BUSER : STD_LOGIC_VECTOR (0 downto 0);
    signal indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter1_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_sig_ioackin_gmem_ARREADY : STD_LOGIC;
    signal ap_pipeline_reg_pp0_iter2_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter3_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter4_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter5_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter6_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter7_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter8_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter9_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter10_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter11_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter12_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter13_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter14_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter15_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter16_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter17_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter18_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter19_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter20_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter21_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter22_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter23_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter24_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter25_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter26_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter27_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter28_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter29_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter30_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter31_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter32_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter33_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter34_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter35_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter36_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter37_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter38_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter39_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter40_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter41_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter42_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter43_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter44_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter45_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter46_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter47_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter48_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter49_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter50_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter51_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter52_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter53_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter54_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter55_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter56_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter57_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter58_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter59_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter60_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter61_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter62_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter63_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter64_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter65_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter66_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter67_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter68_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter69_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter70_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter71_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter72_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter73_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter74_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter75_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter76_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter77_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter78_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter79_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter80_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter81_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter82_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter83_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter84_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter85_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter86_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter87_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter88_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter89_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter90_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter91_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter92_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter93_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter94_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter95_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter96_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter97_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter98_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter99_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter100_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter101_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter102_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter103_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter104_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter105_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter106_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter107_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter108_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter109_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter110_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter111_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter112_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter113_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter114_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter115_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter116_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter117_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter118_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter119_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter120_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter121_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter122_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter123_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter124_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter125_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter126_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter127_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter128_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter129_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter130_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter131_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter132_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter133_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter134_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp0_iter135_indvar_reg_191 : STD_LOGIC_VECTOR (4 downto 0);
    signal indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter1_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter2_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter3_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter4_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter5_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter6_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter7_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter8_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter9_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter10_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter11_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter12_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter13_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter14_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter15_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter16_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter17_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter18_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter19_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter20_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter21_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter22_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter23_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter24_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter25_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter26_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter27_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter28_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter29_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter30_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter31_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter32_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter33_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter34_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter35_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter36_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter37_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter38_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter39_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter40_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter41_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter42_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter43_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter44_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter45_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter46_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter47_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter48_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter49_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter50_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter51_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter52_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter53_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter54_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter55_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter56_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter57_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter58_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter59_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter60_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter61_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter62_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter63_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter64_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter65_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter66_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter67_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter68_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter69_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter70_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter71_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter72_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter73_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter74_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter75_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter76_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter77_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter78_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter79_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter80_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter81_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter82_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter83_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter84_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter85_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter86_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter87_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter88_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter89_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter90_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter91_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter92_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter93_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter94_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter95_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter96_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter97_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter98_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter99_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter100_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter101_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter102_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter103_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter104_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter105_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter106_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter107_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter108_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter109_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter110_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter111_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter112_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter113_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter114_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter115_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter116_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter117_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter118_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter119_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter120_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter121_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter122_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter123_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter124_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter125_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter126_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter127_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter128_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter129_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter130_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter131_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter132_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter133_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter134_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_pipeline_reg_pp1_iter135_indvar7_reg_203 : STD_LOGIC_VECTOR (4 downto 0);
    signal reg_230 : STD_LOGIC_VECTOR (31 downto 0);
    signal global_offset_x_read_reg_435 : STD_LOGIC_VECTOR (31 downto 0);
    signal tmp_fu_234_p1 : STD_LOGIC_VECTOR (5 downto 0);
    signal tmp_reg_440 : STD_LOGIC_VECTOR (5 downto 0);
    signal tmp_1_fu_238_p1 : STD_LOGIC_VECTOR (25 downto 0);
    signal tmp_1_reg_445 : STD_LOGIC_VECTOR (25 downto 0);
    signal tmp_cast_fu_246_p3 : STD_LOGIC_VECTOR (5 downto 0);
    signal tmp_cast_reg_450 : STD_LOGIC_VECTOR (5 downto 0);
    signal arg_x_reg_455 : STD_LOGIC_VECTOR (31 downto 0);
    signal arg_y_reg_461 : STD_LOGIC_VECTOR (31 downto 0);
    signal tmp_6_cast_fu_304_p1 : STD_LOGIC_VECTOR (30 downto 0);
    signal tmp_6_cast_reg_467 : STD_LOGIC_VECTOR (30 downto 0);
    signal exitcond_fu_308_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter1_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter2_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter3_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter4_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter5_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter6_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter7_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter8_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter9_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter10_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter11_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter12_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter13_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter14_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter15_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter16_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter17_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter18_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter19_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter20_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter21_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter22_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter23_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter24_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter25_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter26_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter27_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter28_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter29_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter30_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter31_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter32_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter33_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter34_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter35_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter36_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter37_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter38_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter39_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter40_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter41_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter42_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter43_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter44_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter45_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter46_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter47_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter48_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter49_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter50_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter51_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter52_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter53_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter54_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter55_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter56_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter57_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter58_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter59_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter60_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter61_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter62_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter63_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter64_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter65_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter66_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter67_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter68_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter69_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter70_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter71_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter72_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter73_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter74_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter75_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter76_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter77_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter78_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter79_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter80_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter81_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter82_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter83_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter84_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter85_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter86_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter87_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter88_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter89_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter90_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter91_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter92_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter93_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter94_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter95_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter96_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter97_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter98_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter99_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter100_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter101_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter102_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter103_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter104_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter105_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter106_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter107_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter108_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter109_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter110_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter111_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter112_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter113_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter114_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter115_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter116_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter117_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter118_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter119_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter120_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter121_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter122_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter123_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter124_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter125_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter126_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter127_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter128_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter129_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter130_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter131_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter132_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter133_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp0_iter135_exitcond_reg_472 : STD_LOGIC_VECTOR (0 downto 0);
    signal indvar_next_fu_314_p2 : STD_LOGIC_VECTOR (4 downto 0);
    signal indvar_next_reg_476 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_enable_reg_pp0_iter0 : STD_LOGIC := '0';
    signal isIter0_fu_320_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal exitcond9_fu_336_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter1_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter2_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter3_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter4_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter5_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter6_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter7_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter8_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter9_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter10_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter11_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter12_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter13_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter14_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter15_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter16_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter17_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter18_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter19_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter20_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter21_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter22_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter23_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter24_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter25_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter26_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter27_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter28_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter29_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter30_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter31_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter32_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter33_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter34_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter35_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter36_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter37_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter38_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter39_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter40_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter41_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter42_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter43_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter44_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter45_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter46_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter47_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter48_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter49_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter50_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter51_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter52_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter53_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter54_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter55_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter56_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter57_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter58_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter59_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter60_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter61_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter62_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter63_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter64_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter65_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter66_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter67_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter68_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter69_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter70_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter71_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter72_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter73_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter74_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter75_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter76_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter77_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter78_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter79_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter80_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter81_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter82_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter83_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter84_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter85_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter86_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter87_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter88_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter89_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter90_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter91_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter92_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter93_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter94_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter95_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter96_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter97_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter98_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter99_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter100_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter101_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter102_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter103_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter104_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter105_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter106_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter107_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter108_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter109_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter110_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter111_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter112_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter113_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter114_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter115_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter116_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter117_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter118_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter119_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter120_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter121_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter122_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter123_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter124_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter125_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter126_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter127_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter128_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter129_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter130_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter131_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter132_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter133_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_pipeline_reg_pp1_iter135_exitcond9_reg_485 : STD_LOGIC_VECTOR (0 downto 0);
    signal indvar_next8_fu_342_p2 : STD_LOGIC_VECTOR (4 downto 0);
    signal indvar_next8_reg_489 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_enable_reg_pp1_iter0 : STD_LOGIC := '0';
    signal isIter_fu_348_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal tmp_16_fu_384_p2 : STD_LOGIC_VECTOR (30 downto 0);
    signal tmp_16_reg_498 : STD_LOGIC_VECTOR (30 downto 0);
    signal ap_CS_fsm_state277 : STD_LOGIC_VECTOR (0 downto 0);
    attribute fsm_encoding of ap_CS_fsm_state277 : signal is "none";
    signal ap_sig_ioackin_gmem_AWREADY : STD_LOGIC;
    signal indvar_inc_reg2mem_fu_405_p2 : STD_LOGIC_VECTOR (4 downto 0);
    signal indvar_inc_reg2mem_reg_511 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_CS_fsm_state279 : STD_LOGIC_VECTOR (0 downto 0);
    attribute fsm_encoding of ap_CS_fsm_state279 : signal is "none";
    signal tmp_9_fu_399_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal x0_load_reg_526 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_CS_fsm_state280 : STD_LOGIC_VECTOR (0 downto 0);
    attribute fsm_encoding of ap_CS_fsm_state280 : signal is "none";
    signal y0_load_reg_531 : STD_LOGIC_VECTOR (31 downto 0);
    signal grp_fu_226_p2 : STD_LOGIC_VECTOR (31 downto 0);
    signal tmp_3_reg_536 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_CS_fsm_state284 : STD_LOGIC_VECTOR (0 downto 0);
    attribute fsm_encoding of ap_CS_fsm_state284 : signal is "none";
    signal ap_enable_reg_pp0_iter2 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter3 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter4 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter5 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter6 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter7 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter8 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter9 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter10 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter11 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter12 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter13 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter14 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter15 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter16 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter17 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter18 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter19 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter20 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter21 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter22 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter23 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter24 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter25 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter26 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter27 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter28 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter29 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter30 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter31 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter32 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter33 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter34 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter35 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter36 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter37 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter38 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter39 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter40 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter41 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter42 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter43 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter44 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter45 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter46 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter47 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter48 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter49 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter50 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter51 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter52 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter53 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter54 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter55 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter56 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter57 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter58 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter59 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter60 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter61 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter62 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter63 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter64 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter65 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter66 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter67 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter68 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter69 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter70 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter71 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter72 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter73 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter74 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter75 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter76 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter77 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter78 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter79 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter80 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter81 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter82 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter83 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter84 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter85 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter86 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter87 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter88 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter89 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter90 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter91 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter92 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter93 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter94 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter95 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter96 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter97 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter98 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter99 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter100 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter101 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter102 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter103 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter104 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter105 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter106 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter107 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter108 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter109 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter110 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter111 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter112 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter113 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter114 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter115 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter116 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter117 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter118 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter119 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter120 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter121 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter122 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter123 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter124 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter125 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter126 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter127 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter128 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter129 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter130 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter131 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter132 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter133 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter134 : STD_LOGIC := '0';
    signal ap_enable_reg_pp0_iter136 : STD_LOGIC := '0';
    signal ap_CS_fsm_state139 : STD_LOGIC_VECTOR (0 downto 0);
    attribute fsm_encoding of ap_CS_fsm_state139 : signal is "none";
    signal ap_enable_reg_pp1_iter2 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter3 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter4 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter5 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter6 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter7 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter8 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter9 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter10 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter11 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter12 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter13 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter14 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter15 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter16 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter17 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter18 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter19 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter20 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter21 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter22 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter23 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter24 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter25 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter26 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter27 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter28 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter29 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter30 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter31 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter32 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter33 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter34 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter35 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter36 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter37 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter38 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter39 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter40 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter41 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter42 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter43 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter44 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter45 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter46 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter47 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter48 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter49 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter50 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter51 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter52 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter53 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter54 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter55 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter56 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter57 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter58 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter59 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter60 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter61 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter62 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter63 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter64 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter65 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter66 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter67 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter68 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter69 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter70 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter71 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter72 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter73 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter74 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter75 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter76 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter77 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter78 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter79 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter80 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter81 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter82 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter83 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter84 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter85 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter86 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter87 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter88 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter89 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter90 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter91 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter92 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter93 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter94 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter95 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter96 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter97 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter98 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter99 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter100 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter101 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter102 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter103 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter104 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter105 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter106 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter107 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter108 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter109 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter110 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter111 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter112 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter113 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter114 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter115 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter116 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter117 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter118 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter119 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter120 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter121 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter122 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter123 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter124 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter125 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter126 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter127 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter128 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter129 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter130 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter131 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter132 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter133 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter134 : STD_LOGIC := '0';
    signal ap_enable_reg_pp1_iter136 : STD_LOGIC := '0';
    signal indvar_phi_fu_195_p4 : STD_LOGIC_VECTOR (4 downto 0);
    signal indvar7_phi_fu_207_p4 : STD_LOGIC_VECTOR (4 downto 0);
    signal indvar_reg2mem44_0_i_reg_215 : STD_LOGIC_VECTOR (4 downto 0);
    signal ap_sig_ioackin_gmem_WREADY : STD_LOGIC;
    signal indvar_cast_fu_326_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal indvar7_cast_fu_354_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal tmp_2_cast1_fu_425_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal tmp_10_fu_264_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal tmp_11_fu_284_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal tmp_17_fu_389_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_reg_ioackin_gmem_ARREADY : STD_LOGIC := '0';
    signal ap_reg_ioackin_gmem_AWREADY : STD_LOGIC := '0';
    signal ap_reg_ioackin_gmem_WREADY : STD_LOGIC := '0';
    signal ap_CS_fsm_state281 : STD_LOGIC_VECTOR (0 downto 0);
    attribute fsm_encoding of ap_CS_fsm_state281 : signal is "none";
    signal tmp_6_fu_242_p1 : STD_LOGIC_VECTOR (1 downto 0);
    signal tmp_4_fu_254_p4 : STD_LOGIC_VECTOR (29 downto 0);
    signal tmp_5_fu_274_p4 : STD_LOGIC_VECTOR (29 downto 0);
    signal tmp_12_fu_294_p4 : STD_LOGIC_VECTOR (29 downto 0);
    signal tmp_7_fu_364_p3 : STD_LOGIC_VECTOR (29 downto 0);
    signal tmp_13_fu_371_p1 : STD_LOGIC_VECTOR (29 downto 0);
    signal tmp_14_fu_374_p2 : STD_LOGIC_VECTOR (29 downto 0);
    signal tmp_15_fu_380_p1 : STD_LOGIC_VECTOR (30 downto 0);
    signal indvar_reg2mem44_0_i_1_fu_411_p1 : STD_LOGIC_VECTOR (5 downto 0);
    signal tmp1_fu_415_p2 : STD_LOGIC_VECTOR (5 downto 0);
    signal tmp_2_fu_420_p2 : STD_LOGIC_VECTOR (5 downto 0);
    signal ap_NS_fsm : STD_LOGIC_VECTOR (143 downto 0);
    signal ap_condition_1658 : BOOLEAN;
    signal ap_condition_1670 : BOOLEAN;

    component gpu_fadd_32ns_32nbkb IS
    generic (
        ID : INTEGER;
        NUM_STAGE : INTEGER;
        din0_WIDTH : INTEGER;
        din1_WIDTH : INTEGER;
        dout_WIDTH : INTEGER );
    port (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        din0 : IN STD_LOGIC_VECTOR (31 downto 0);
        din1 : IN STD_LOGIC_VECTOR (31 downto 0);
        ce : IN STD_LOGIC;
        dout : OUT STD_LOGIC_VECTOR (31 downto 0) );
    end component;


    component gpu_x0 IS
    generic (
        DataWidth : INTEGER;
        AddressRange : INTEGER;
        AddressWidth : INTEGER );
    port (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        address0 : IN STD_LOGIC_VECTOR (3 downto 0);
        ce0 : IN STD_LOGIC;
        we0 : IN STD_LOGIC;
        d0 : IN STD_LOGIC_VECTOR (31 downto 0);
        q0 : OUT STD_LOGIC_VECTOR (31 downto 0) );
    end component;


    component gpu_control_s_axi IS
    generic (
        C_S_AXI_ADDR_WIDTH : INTEGER;
        C_S_AXI_DATA_WIDTH : INTEGER );
    port (
        AWVALID : IN STD_LOGIC;
        AWREADY : OUT STD_LOGIC;
        AWADDR : IN STD_LOGIC_VECTOR (C_S_AXI_ADDR_WIDTH-1 downto 0);
        WVALID : IN STD_LOGIC;
        WREADY : OUT STD_LOGIC;
        WDATA : IN STD_LOGIC_VECTOR (C_S_AXI_DATA_WIDTH-1 downto 0);
        WSTRB : IN STD_LOGIC_VECTOR (C_S_AXI_DATA_WIDTH/8-1 downto 0);
        ARVALID : IN STD_LOGIC;
        ARREADY : OUT STD_LOGIC;
        ARADDR : IN STD_LOGIC_VECTOR (C_S_AXI_ADDR_WIDTH-1 downto 0);
        RVALID : OUT STD_LOGIC;
        RREADY : IN STD_LOGIC;
        RDATA : OUT STD_LOGIC_VECTOR (C_S_AXI_DATA_WIDTH-1 downto 0);
        RRESP : OUT STD_LOGIC_VECTOR (1 downto 0);
        BVALID : OUT STD_LOGIC;
        BREADY : IN STD_LOGIC;
        BRESP : OUT STD_LOGIC_VECTOR (1 downto 0);
        ACLK : IN STD_LOGIC;
        ARESET : IN STD_LOGIC;
        ACLK_EN : IN STD_LOGIC;
        ap_start : OUT STD_LOGIC;
        interrupt : OUT STD_LOGIC;
        ap_ready : IN STD_LOGIC;
        ap_done : IN STD_LOGIC;
        ap_idle : IN STD_LOGIC;
        group_id_x : OUT STD_LOGIC_VECTOR (31 downto 0);
        group_id_y : OUT STD_LOGIC_VECTOR (31 downto 0);
        group_id_z : OUT STD_LOGIC_VECTOR (31 downto 0);
        global_offset_x : OUT STD_LOGIC_VECTOR (31 downto 0);
        global_offset_y : OUT STD_LOGIC_VECTOR (31 downto 0);
        global_offset_z : OUT STD_LOGIC_VECTOR (31 downto 0);
        x : OUT STD_LOGIC_VECTOR (31 downto 0);
        y : OUT STD_LOGIC_VECTOR (31 downto 0);
        z : OUT STD_LOGIC_VECTOR (31 downto 0) );
    end component;


    component gpu_gmem_m_axi IS
    generic (
        USER_DW : INTEGER;
        USER_AW : INTEGER;
        USER_MAXREQS : INTEGER;
        NUM_READ_OUTSTANDING : INTEGER;
        NUM_WRITE_OUTSTANDING : INTEGER;
        MAX_READ_BURST_LENGTH : INTEGER;
        MAX_WRITE_BURST_LENGTH : INTEGER;
        C_M_AXI_ID_WIDTH : INTEGER;
        C_M_AXI_ADDR_WIDTH : INTEGER;
        C_M_AXI_DATA_WIDTH : INTEGER;
        C_M_AXI_AWUSER_WIDTH : INTEGER;
        C_M_AXI_ARUSER_WIDTH : INTEGER;
        C_M_AXI_WUSER_WIDTH : INTEGER;
        C_M_AXI_RUSER_WIDTH : INTEGER;
        C_M_AXI_BUSER_WIDTH : INTEGER;
        C_TARGET_ADDR : INTEGER;
        C_USER_VALUE : INTEGER;
        C_PROT_VALUE : INTEGER;
        C_CACHE_VALUE : INTEGER );
    port (
        AWVALID : OUT STD_LOGIC;
        AWREADY : IN STD_LOGIC;
        AWADDR : OUT STD_LOGIC_VECTOR (C_M_AXI_ADDR_WIDTH-1 downto 0);
        AWID : OUT STD_LOGIC_VECTOR (C_M_AXI_ID_WIDTH-1 downto 0);
        AWLEN : OUT STD_LOGIC_VECTOR (7 downto 0);
        AWSIZE : OUT STD_LOGIC_VECTOR (2 downto 0);
        AWBURST : OUT STD_LOGIC_VECTOR (1 downto 0);
        AWLOCK : OUT STD_LOGIC_VECTOR (1 downto 0);
        AWCACHE : OUT STD_LOGIC_VECTOR (3 downto 0);
        AWPROT : OUT STD_LOGIC_VECTOR (2 downto 0);
        AWQOS : OUT STD_LOGIC_VECTOR (3 downto 0);
        AWREGION : OUT STD_LOGIC_VECTOR (3 downto 0);
        AWUSER : OUT STD_LOGIC_VECTOR (C_M_AXI_AWUSER_WIDTH-1 downto 0);
        WVALID : OUT STD_LOGIC;
        WREADY : IN STD_LOGIC;
        WDATA : OUT STD_LOGIC_VECTOR (C_M_AXI_DATA_WIDTH-1 downto 0);
        WSTRB : OUT STD_LOGIC_VECTOR (C_M_AXI_DATA_WIDTH/8-1 downto 0);
        WLAST : OUT STD_LOGIC;
        WID : OUT STD_LOGIC_VECTOR (C_M_AXI_ID_WIDTH-1 downto 0);
        WUSER : OUT STD_LOGIC_VECTOR (C_M_AXI_WUSER_WIDTH-1 downto 0);
        ARVALID : OUT STD_LOGIC;
        ARREADY : IN STD_LOGIC;
        ARADDR : OUT STD_LOGIC_VECTOR (C_M_AXI_ADDR_WIDTH-1 downto 0);
        ARID : OUT STD_LOGIC_VECTOR (C_M_AXI_ID_WIDTH-1 downto 0);
        ARLEN : OUT STD_LOGIC_VECTOR (7 downto 0);
        ARSIZE : OUT STD_LOGIC_VECTOR (2 downto 0);
        ARBURST : OUT STD_LOGIC_VECTOR (1 downto 0);
        ARLOCK : OUT STD_LOGIC_VECTOR (1 downto 0);
        ARCACHE : OUT STD_LOGIC_VECTOR (3 downto 0);
        ARPROT : OUT STD_LOGIC_VECTOR (2 downto 0);
        ARQOS : OUT STD_LOGIC_VECTOR (3 downto 0);
        ARREGION : OUT STD_LOGIC_VECTOR (3 downto 0);
        ARUSER : OUT STD_LOGIC_VECTOR (C_M_AXI_ARUSER_WIDTH-1 downto 0);
        RVALID : IN STD_LOGIC;
        RREADY : OUT STD_LOGIC;
        RDATA : IN STD_LOGIC_VECTOR (C_M_AXI_DATA_WIDTH-1 downto 0);
        RLAST : IN STD_LOGIC;
        RID : IN STD_LOGIC_VECTOR (C_M_AXI_ID_WIDTH-1 downto 0);
        RUSER : IN STD_LOGIC_VECTOR (C_M_AXI_RUSER_WIDTH-1 downto 0);
        RRESP : IN STD_LOGIC_VECTOR (1 downto 0);
        BVALID : IN STD_LOGIC;
        BREADY : OUT STD_LOGIC;
        BRESP : IN STD_LOGIC_VECTOR (1 downto 0);
        BID : IN STD_LOGIC_VECTOR (C_M_AXI_ID_WIDTH-1 downto 0);
        BUSER : IN STD_LOGIC_VECTOR (C_M_AXI_BUSER_WIDTH-1 downto 0);
        ACLK : IN STD_LOGIC;
        ARESET : IN STD_LOGIC;
        ACLK_EN : IN STD_LOGIC;
        I_ARVALID : IN STD_LOGIC;
        I_ARREADY : OUT STD_LOGIC;
        I_ARADDR : IN STD_LOGIC_VECTOR (31 downto 0);
        I_ARID : IN STD_LOGIC_VECTOR (0 downto 0);
        I_ARLEN : IN STD_LOGIC_VECTOR (31 downto 0);
        I_ARSIZE : IN STD_LOGIC_VECTOR (2 downto 0);
        I_ARLOCK : IN STD_LOGIC_VECTOR (1 downto 0);
        I_ARCACHE : IN STD_LOGIC_VECTOR (3 downto 0);
        I_ARQOS : IN STD_LOGIC_VECTOR (3 downto 0);
        I_ARPROT : IN STD_LOGIC_VECTOR (2 downto 0);
        I_ARUSER : IN STD_LOGIC_VECTOR (0 downto 0);
        I_ARBURST : IN STD_LOGIC_VECTOR (1 downto 0);
        I_ARREGION : IN STD_LOGIC_VECTOR (3 downto 0);
        I_RVALID : OUT STD_LOGIC;
        I_RREADY : IN STD_LOGIC;
        I_RDATA : OUT STD_LOGIC_VECTOR (31 downto 0);
        I_RID : OUT STD_LOGIC_VECTOR (0 downto 0);
        I_RUSER : OUT STD_LOGIC_VECTOR (0 downto 0);
        I_RRESP : OUT STD_LOGIC_VECTOR (1 downto 0);
        I_RLAST : OUT STD_LOGIC;
        I_AWVALID : IN STD_LOGIC;
        I_AWREADY : OUT STD_LOGIC;
        I_AWADDR : IN STD_LOGIC_VECTOR (31 downto 0);
        I_AWID : IN STD_LOGIC_VECTOR (0 downto 0);
        I_AWLEN : IN STD_LOGIC_VECTOR (31 downto 0);
        I_AWSIZE : IN STD_LOGIC_VECTOR (2 downto 0);
        I_AWLOCK : IN STD_LOGIC_VECTOR (1 downto 0);
        I_AWCACHE : IN STD_LOGIC_VECTOR (3 downto 0);
        I_AWQOS : IN STD_LOGIC_VECTOR (3 downto 0);
        I_AWPROT : IN STD_LOGIC_VECTOR (2 downto 0);
        I_AWUSER : IN STD_LOGIC_VECTOR (0 downto 0);
        I_AWBURST : IN STD_LOGIC_VECTOR (1 downto 0);
        I_AWREGION : IN STD_LOGIC_VECTOR (3 downto 0);
        I_WVALID : IN STD_LOGIC;
        I_WREADY : OUT STD_LOGIC;
        I_WDATA : IN STD_LOGIC_VECTOR (31 downto 0);
        I_WID : IN STD_LOGIC_VECTOR (0 downto 0);
        I_WUSER : IN STD_LOGIC_VECTOR (0 downto 0);
        I_WLAST : IN STD_LOGIC;
        I_WSTRB : IN STD_LOGIC_VECTOR (3 downto 0);
        I_BVALID : OUT STD_LOGIC;
        I_BREADY : IN STD_LOGIC;
        I_BRESP : OUT STD_LOGIC_VECTOR (1 downto 0);
        I_BID : OUT STD_LOGIC_VECTOR (0 downto 0);
        I_BUSER : OUT STD_LOGIC_VECTOR (0 downto 0) );
    end component;



begin
    x0_U : component gpu_x0
    generic map (
        DataWidth => 32,
        AddressRange => 16,
        AddressWidth => 4)
    port map (
        clk => ap_clk,
        reset => ap_rst_n_inv,
        address0 => x0_address0,
        ce0 => x0_ce0,
        we0 => x0_we0,
        d0 => x0_d0,
        q0 => x0_q0);

    y0_U : component gpu_x0
    generic map (
        DataWidth => 32,
        AddressRange => 16,
        AddressWidth => 4)
    port map (
        clk => ap_clk,
        reset => ap_rst_n_inv,
        address0 => y0_address0,
        ce0 => y0_ce0,
        we0 => y0_we0,
        d0 => y0_d0,
        q0 => y0_q0);

    gpu_control_s_axi_U : component gpu_control_s_axi
    generic map (
        C_S_AXI_ADDR_WIDTH => C_S_AXI_CONTROL_ADDR_WIDTH,
        C_S_AXI_DATA_WIDTH => C_S_AXI_CONTROL_DATA_WIDTH)
    port map (
        AWVALID => s_axi_control_AWVALID,
        AWREADY => s_axi_control_AWREADY,
        AWADDR => s_axi_control_AWADDR,
        WVALID => s_axi_control_WVALID,
        WREADY => s_axi_control_WREADY,
        WDATA => s_axi_control_WDATA,
        WSTRB => s_axi_control_WSTRB,
        ARVALID => s_axi_control_ARVALID,
        ARREADY => s_axi_control_ARREADY,
        ARADDR => s_axi_control_ARADDR,
        RVALID => s_axi_control_RVALID,
        RREADY => s_axi_control_RREADY,
        RDATA => s_axi_control_RDATA,
        RRESP => s_axi_control_RRESP,
        BVALID => s_axi_control_BVALID,
        BREADY => s_axi_control_BREADY,
        BRESP => s_axi_control_BRESP,
        ACLK => ap_clk,
        ARESET => ap_rst_n_inv,
        ACLK_EN => ap_const_logic_1,
        ap_start => ap_start,
        interrupt => interrupt,
        ap_ready => ap_ready,
        ap_done => ap_done,
        ap_idle => ap_idle,
        group_id_x => group_id_x,
        group_id_y => group_id_y,
        group_id_z => group_id_z,
        global_offset_x => global_offset_x,
        global_offset_y => global_offset_y,
        global_offset_z => global_offset_z,
        x => x,
        y => y,
        z => z);

    gpu_gmem_m_axi_U : component gpu_gmem_m_axi
    generic map (
        USER_DW => 32,
        USER_AW => 32,
        USER_MAXREQS => 133,
        NUM_READ_OUTSTANDING => 16,
        NUM_WRITE_OUTSTANDING => 16,
        MAX_READ_BURST_LENGTH => 16,
        MAX_WRITE_BURST_LENGTH => 16,
        C_M_AXI_ID_WIDTH => C_M_AXI_GMEM_ID_WIDTH,
        C_M_AXI_ADDR_WIDTH => C_M_AXI_GMEM_ADDR_WIDTH,
        C_M_AXI_DATA_WIDTH => C_M_AXI_GMEM_DATA_WIDTH,
        C_M_AXI_AWUSER_WIDTH => C_M_AXI_GMEM_AWUSER_WIDTH,
        C_M_AXI_ARUSER_WIDTH => C_M_AXI_GMEM_ARUSER_WIDTH,
        C_M_AXI_WUSER_WIDTH => C_M_AXI_GMEM_WUSER_WIDTH,
        C_M_AXI_RUSER_WIDTH => C_M_AXI_GMEM_RUSER_WIDTH,
        C_M_AXI_BUSER_WIDTH => C_M_AXI_GMEM_BUSER_WIDTH,
        C_TARGET_ADDR => C_M_AXI_GMEM_TARGET_ADDR,
        C_USER_VALUE => C_M_AXI_GMEM_USER_VALUE,
        C_PROT_VALUE => C_M_AXI_GMEM_PROT_VALUE,
        C_CACHE_VALUE => C_M_AXI_GMEM_CACHE_VALUE)
    port map (
        AWVALID => m_axi_gmem_AWVALID,
        AWREADY => m_axi_gmem_AWREADY,
        AWADDR => m_axi_gmem_AWADDR,
        AWID => m_axi_gmem_AWID,
        AWLEN => m_axi_gmem_AWLEN,
        AWSIZE => m_axi_gmem_AWSIZE,
        AWBURST => m_axi_gmem_AWBURST,
        AWLOCK => m_axi_gmem_AWLOCK,
        AWCACHE => m_axi_gmem_AWCACHE,
        AWPROT => m_axi_gmem_AWPROT,
        AWQOS => m_axi_gmem_AWQOS,
        AWREGION => m_axi_gmem_AWREGION,
        AWUSER => m_axi_gmem_AWUSER,
        WVALID => m_axi_gmem_WVALID,
        WREADY => m_axi_gmem_WREADY,
        WDATA => m_axi_gmem_WDATA,
        WSTRB => m_axi_gmem_WSTRB,
        WLAST => m_axi_gmem_WLAST,
        WID => m_axi_gmem_WID,
        WUSER => m_axi_gmem_WUSER,
        ARVALID => m_axi_gmem_ARVALID,
        ARREADY => m_axi_gmem_ARREADY,
        ARADDR => m_axi_gmem_ARADDR,
        ARID => m_axi_gmem_ARID,
        ARLEN => m_axi_gmem_ARLEN,
        ARSIZE => m_axi_gmem_ARSIZE,
        ARBURST => m_axi_gmem_ARBURST,
        ARLOCK => m_axi_gmem_ARLOCK,
        ARCACHE => m_axi_gmem_ARCACHE,
        ARPROT => m_axi_gmem_ARPROT,
        ARQOS => m_axi_gmem_ARQOS,
        ARREGION => m_axi_gmem_ARREGION,
        ARUSER => m_axi_gmem_ARUSER,
        RVALID => m_axi_gmem_RVALID,
        RREADY => m_axi_gmem_RREADY,
        RDATA => m_axi_gmem_RDATA,
        RLAST => m_axi_gmem_RLAST,
        RID => m_axi_gmem_RID,
        RUSER => m_axi_gmem_RUSER,
        RRESP => m_axi_gmem_RRESP,
        BVALID => m_axi_gmem_BVALID,
        BREADY => m_axi_gmem_BREADY,
        BRESP => m_axi_gmem_BRESP,
        BID => m_axi_gmem_BID,
        BUSER => m_axi_gmem_BUSER,
        ACLK => ap_clk,
        ARESET => ap_rst_n_inv,
        ACLK_EN => ap_const_logic_1,
        I_ARVALID => gmem_ARVALID,
        I_ARREADY => gmem_ARREADY,
        I_ARADDR => gmem_ARADDR,
        I_ARID => ap_const_lv1_0,
        I_ARLEN => ap_const_lv32_10,
        I_ARSIZE => ap_const_lv3_0,
        I_ARLOCK => ap_const_lv2_0,
        I_ARCACHE => ap_const_lv4_0,
        I_ARQOS => ap_const_lv4_0,
        I_ARPROT => ap_const_lv3_0,
        I_ARUSER => ap_const_lv1_0,
        I_ARBURST => ap_const_lv2_0,
        I_ARREGION => ap_const_lv4_0,
        I_RVALID => gmem_RVALID,
        I_RREADY => gmem_RREADY,
        I_RDATA => gmem_RDATA,
        I_RID => gmem_RID,
        I_RUSER => gmem_RUSER,
        I_RRESP => gmem_RRESP,
        I_RLAST => gmem_RLAST,
        I_AWVALID => gmem_AWVALID,
        I_AWREADY => gmem_AWREADY,
        I_AWADDR => tmp_17_fu_389_p1,
        I_AWID => ap_const_lv1_0,
        I_AWLEN => ap_const_lv32_10,
        I_AWSIZE => ap_const_lv3_0,
        I_AWLOCK => ap_const_lv2_0,
        I_AWCACHE => ap_const_lv4_0,
        I_AWQOS => ap_const_lv4_0,
        I_AWPROT => ap_const_lv3_0,
        I_AWUSER => ap_const_lv1_0,
        I_AWBURST => ap_const_lv2_0,
        I_AWREGION => ap_const_lv4_0,
        I_WVALID => gmem_WVALID,
        I_WREADY => gmem_WREADY,
        I_WDATA => gmem_WDATA,
        I_WID => ap_const_lv1_0,
        I_WUSER => ap_const_lv1_0,
        I_WLAST => ap_const_logic_0,
        I_WSTRB => ap_const_lv4_F,
        I_BVALID => gmem_BVALID,
        I_BREADY => gmem_BREADY,
        I_BRESP => gmem_BRESP,
        I_BID => gmem_BID,
        I_BUSER => gmem_BUSER);

    gpu_fadd_32ns_32nbkb_U1 : component gpu_fadd_32ns_32nbkb
    generic map (
        ID => 1,
        NUM_STAGE => 4,
        din0_WIDTH => 32,
        din1_WIDTH => 32,
        dout_WIDTH => 32)
    port map (
        clk => ap_clk,
        reset => ap_rst_n_inv,
        din0 => x0_load_reg_526,
        din1 => y0_load_reg_531,
        ce => ap_const_logic_1,
        dout => grp_fu_226_p2);





    ap_CS_fsm_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_CS_fsm <= ap_ST_fsm_state1;
            else
                ap_CS_fsm <= ap_NS_fsm;
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter0_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter0 <= ap_const_logic_0;
            else
                if (((ap_const_lv1_1 = ap_CS_fsm_pp0_stage0) and not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))) and not((ap_const_lv1_0 = exitcond_fu_308_p2)))) then 
                    ap_enable_reg_pp0_iter0 <= ap_const_logic_0;
                elsif (((ap_CS_fsm_state1 = ap_const_lv1_1) and not((ap_start = ap_const_logic_0)))) then 
                    ap_enable_reg_pp0_iter0 <= ap_const_logic_1;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter1_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter1 <= ap_const_logic_0;
            else
                if (((ap_const_lv1_1 = ap_CS_fsm_pp0_stage0) and not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_lv1_0 = exitcond_fu_308_p2))) then 
                    ap_enable_reg_pp0_iter1 <= ap_const_logic_1;
                elsif ((((ap_CS_fsm_state1 = ap_const_lv1_1) and not((ap_start = ap_const_logic_0))) or ((ap_const_lv1_1 = ap_CS_fsm_pp0_stage0) and not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))) and not((ap_const_lv1_0 = exitcond_fu_308_p2))))) then 
                    ap_enable_reg_pp0_iter1 <= ap_const_logic_0;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter10_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter10 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter100_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter100 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter100 <= ap_enable_reg_pp0_iter99;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter101_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter101 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter101 <= ap_enable_reg_pp0_iter100;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter102_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter102 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter102 <= ap_enable_reg_pp0_iter101;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter103_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter103 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter103 <= ap_enable_reg_pp0_iter102;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter104_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter104 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter104 <= ap_enable_reg_pp0_iter103;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter105_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter105 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter105 <= ap_enable_reg_pp0_iter104;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter106_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter106 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter106 <= ap_enable_reg_pp0_iter105;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter107_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter107 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter107 <= ap_enable_reg_pp0_iter106;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter108_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter108 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter108 <= ap_enable_reg_pp0_iter107;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter109_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter109 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter109 <= ap_enable_reg_pp0_iter108;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter11_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter11 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter110_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter110 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter110 <= ap_enable_reg_pp0_iter109;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter111_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter111 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter111 <= ap_enable_reg_pp0_iter110;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter112_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter112 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter112 <= ap_enable_reg_pp0_iter111;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter113_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter113 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter113 <= ap_enable_reg_pp0_iter112;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter114_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter114 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter114 <= ap_enable_reg_pp0_iter113;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter115_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter115 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter115 <= ap_enable_reg_pp0_iter114;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter116_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter116 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter116 <= ap_enable_reg_pp0_iter115;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter117_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter117 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter117 <= ap_enable_reg_pp0_iter116;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter118_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter118 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter118 <= ap_enable_reg_pp0_iter117;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter119_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter119 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter119 <= ap_enable_reg_pp0_iter118;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter12_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter12 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter120_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter120 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter120 <= ap_enable_reg_pp0_iter119;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter121_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter121 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter121 <= ap_enable_reg_pp0_iter120;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter122_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter122 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter122 <= ap_enable_reg_pp0_iter121;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter123_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter123 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter123 <= ap_enable_reg_pp0_iter122;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter124_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter124 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter124 <= ap_enable_reg_pp0_iter123;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter125_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter125 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter125 <= ap_enable_reg_pp0_iter124;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter126_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter126 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter126 <= ap_enable_reg_pp0_iter125;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter127_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter127 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter127 <= ap_enable_reg_pp0_iter126;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter128_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter128 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter128 <= ap_enable_reg_pp0_iter127;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter129_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter129 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter129 <= ap_enable_reg_pp0_iter128;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter13_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter13 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter130_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter130 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter130 <= ap_enable_reg_pp0_iter129;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter131_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter131 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter131 <= ap_enable_reg_pp0_iter130;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter132_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter132 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter132 <= ap_enable_reg_pp0_iter131;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter133_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter133 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter133 <= ap_enable_reg_pp0_iter132;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter134_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter134 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter134 <= ap_enable_reg_pp0_iter133;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter135_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter135 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter135 <= ap_enable_reg_pp0_iter134;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter136_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter136 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter136 <= ap_enable_reg_pp0_iter135;
                elsif (((ap_CS_fsm_state1 = ap_const_lv1_1) and not((ap_start = ap_const_logic_0)))) then 
                    ap_enable_reg_pp0_iter136 <= ap_const_logic_0;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter14_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter14 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter15_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter15 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter16_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter16 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter17_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter17 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter18_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter18 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter19_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter19 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter2_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter2 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter20_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter20 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter21_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter21 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter22_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter22 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter23_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter23 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter23 <= ap_enable_reg_pp0_iter22;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter24_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter24 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter24 <= ap_enable_reg_pp0_iter23;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter25_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter25 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter25 <= ap_enable_reg_pp0_iter24;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter26_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter26 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter26 <= ap_enable_reg_pp0_iter25;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter27_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter27 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter27 <= ap_enable_reg_pp0_iter26;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter28_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter28 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter28 <= ap_enable_reg_pp0_iter27;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter29_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter29 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter29 <= ap_enable_reg_pp0_iter28;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter3_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter3 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter30_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter30 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter30 <= ap_enable_reg_pp0_iter29;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter31_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter31 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter31 <= ap_enable_reg_pp0_iter30;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter32_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter32 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter32 <= ap_enable_reg_pp0_iter31;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter33_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter33 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter33 <= ap_enable_reg_pp0_iter32;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter34_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter34 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter34 <= ap_enable_reg_pp0_iter33;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter35_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter35 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter35 <= ap_enable_reg_pp0_iter34;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter36_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter36 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter36 <= ap_enable_reg_pp0_iter35;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter37_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter37 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter37 <= ap_enable_reg_pp0_iter36;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter38_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter38 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter38 <= ap_enable_reg_pp0_iter37;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter39_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter39 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter39 <= ap_enable_reg_pp0_iter38;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter4_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter4 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter40_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter40 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter40 <= ap_enable_reg_pp0_iter39;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter41_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter41 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter41 <= ap_enable_reg_pp0_iter40;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter42_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter42 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter42 <= ap_enable_reg_pp0_iter41;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter43_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter43 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter43 <= ap_enable_reg_pp0_iter42;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter44_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter44 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter44 <= ap_enable_reg_pp0_iter43;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter45_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter45 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter45 <= ap_enable_reg_pp0_iter44;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter46_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter46 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter46 <= ap_enable_reg_pp0_iter45;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter47_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter47 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter47 <= ap_enable_reg_pp0_iter46;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter48_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter48 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter48 <= ap_enable_reg_pp0_iter47;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter49_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter49 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter49 <= ap_enable_reg_pp0_iter48;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter5_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter5 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter50_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter50 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter50 <= ap_enable_reg_pp0_iter49;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter51_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter51 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter51 <= ap_enable_reg_pp0_iter50;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter52_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter52 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter52 <= ap_enable_reg_pp0_iter51;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter53_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter53 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter53 <= ap_enable_reg_pp0_iter52;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter54_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter54 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter54 <= ap_enable_reg_pp0_iter53;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter55_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter55 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter55 <= ap_enable_reg_pp0_iter54;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter56_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter56 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter56 <= ap_enable_reg_pp0_iter55;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter57_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter57 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter57 <= ap_enable_reg_pp0_iter56;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter58_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter58 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter58 <= ap_enable_reg_pp0_iter57;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter59_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter59 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter59 <= ap_enable_reg_pp0_iter58;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter6_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter6 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter60_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter60 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter60 <= ap_enable_reg_pp0_iter59;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter61_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter61 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter61 <= ap_enable_reg_pp0_iter60;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter62_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter62 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter62 <= ap_enable_reg_pp0_iter61;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter63_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter63 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter63 <= ap_enable_reg_pp0_iter62;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter64_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter64 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter64 <= ap_enable_reg_pp0_iter63;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter65_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter65 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter65 <= ap_enable_reg_pp0_iter64;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter66_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter66 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter66 <= ap_enable_reg_pp0_iter65;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter67_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter67 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter67 <= ap_enable_reg_pp0_iter66;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter68_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter68 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter68 <= ap_enable_reg_pp0_iter67;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter69_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter69 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter69 <= ap_enable_reg_pp0_iter68;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter7_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter7 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter70_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter70 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter70 <= ap_enable_reg_pp0_iter69;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter71_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter71 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter71 <= ap_enable_reg_pp0_iter70;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter72_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter72 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter72 <= ap_enable_reg_pp0_iter71;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter73_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter73 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter73 <= ap_enable_reg_pp0_iter72;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter74_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter74 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter74 <= ap_enable_reg_pp0_iter73;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter75_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter75 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter75 <= ap_enable_reg_pp0_iter74;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter76_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter76 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter76 <= ap_enable_reg_pp0_iter75;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter77_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter77 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter77 <= ap_enable_reg_pp0_iter76;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter78_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter78 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter78 <= ap_enable_reg_pp0_iter77;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter79_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter79 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter79 <= ap_enable_reg_pp0_iter78;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter8_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter8 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter80_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter80 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter80 <= ap_enable_reg_pp0_iter79;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter81_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter81 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter81 <= ap_enable_reg_pp0_iter80;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter82_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter82 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter82 <= ap_enable_reg_pp0_iter81;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter83_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter83 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter83 <= ap_enable_reg_pp0_iter82;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter84_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter84 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter84 <= ap_enable_reg_pp0_iter83;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter85_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter85 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter85 <= ap_enable_reg_pp0_iter84;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter86_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter86 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter86 <= ap_enable_reg_pp0_iter85;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter87_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter87 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter87 <= ap_enable_reg_pp0_iter86;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter88_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter88 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter88 <= ap_enable_reg_pp0_iter87;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter89_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter89 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter89 <= ap_enable_reg_pp0_iter88;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter9_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter9 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter90_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter90 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter90 <= ap_enable_reg_pp0_iter89;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter91_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter91 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter91 <= ap_enable_reg_pp0_iter90;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter92_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter92 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter92 <= ap_enable_reg_pp0_iter91;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter93_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter93 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter93 <= ap_enable_reg_pp0_iter92;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter94_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter94 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter94 <= ap_enable_reg_pp0_iter93;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter95_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter95 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter95 <= ap_enable_reg_pp0_iter94;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter96_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter96 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter96 <= ap_enable_reg_pp0_iter95;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter97_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter97 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter97 <= ap_enable_reg_pp0_iter96;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter98_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter98 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter98 <= ap_enable_reg_pp0_iter97;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter99_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter99 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp0_iter99 <= ap_enable_reg_pp0_iter98;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter0_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter0 <= ap_const_logic_0;
            else
                if (((ap_const_lv1_1 = ap_CS_fsm_pp1_stage0) and not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))) and not((ap_const_lv1_0 = exitcond9_fu_336_p2)))) then 
                    ap_enable_reg_pp1_iter0 <= ap_const_logic_0;
                elsif (((ap_const_lv1_1 = ap_CS_fsm_state139))) then 
                    ap_enable_reg_pp1_iter0 <= ap_const_logic_1;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter1_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter1 <= ap_const_logic_0;
            else
                if (((ap_const_lv1_1 = ap_CS_fsm_pp1_stage0) and not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_lv1_0 = exitcond9_fu_336_p2))) then 
                    ap_enable_reg_pp1_iter1 <= ap_const_logic_1;
                elsif ((((ap_const_lv1_1 = ap_CS_fsm_state139)) or ((ap_const_lv1_1 = ap_CS_fsm_pp1_stage0) and not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))) and not((ap_const_lv1_0 = exitcond9_fu_336_p2))))) then 
                    ap_enable_reg_pp1_iter1 <= ap_const_logic_0;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter10_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter10 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter10 <= ap_enable_reg_pp1_iter9;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter100_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter100 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter100 <= ap_enable_reg_pp1_iter99;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter101_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter101 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter101 <= ap_enable_reg_pp1_iter100;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter102_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter102 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter102 <= ap_enable_reg_pp1_iter101;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter103_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter103 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter103 <= ap_enable_reg_pp1_iter102;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter104_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter104 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter104 <= ap_enable_reg_pp1_iter103;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter105_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter105 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter105 <= ap_enable_reg_pp1_iter104;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter106_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter106 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter106 <= ap_enable_reg_pp1_iter105;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter107_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter107 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter107 <= ap_enable_reg_pp1_iter106;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter108_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter108 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter108 <= ap_enable_reg_pp1_iter107;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter109_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter109 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter109 <= ap_enable_reg_pp1_iter108;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter11_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter11 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter11 <= ap_enable_reg_pp1_iter10;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter110_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter110 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter110 <= ap_enable_reg_pp1_iter109;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter111_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter111 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter111 <= ap_enable_reg_pp1_iter110;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter112_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter112 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter112 <= ap_enable_reg_pp1_iter111;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter113_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter113 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter113 <= ap_enable_reg_pp1_iter112;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter114_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter114 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter114 <= ap_enable_reg_pp1_iter113;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter115_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter115 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter115 <= ap_enable_reg_pp1_iter114;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter116_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter116 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter116 <= ap_enable_reg_pp1_iter115;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter117_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter117 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter117 <= ap_enable_reg_pp1_iter116;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter118_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter118 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter118 <= ap_enable_reg_pp1_iter117;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter119_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter119 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter119 <= ap_enable_reg_pp1_iter118;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter12_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter12 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter12 <= ap_enable_reg_pp1_iter11;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter120_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter120 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter120 <= ap_enable_reg_pp1_iter119;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter121_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter121 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter121 <= ap_enable_reg_pp1_iter120;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter122_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter122 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter122 <= ap_enable_reg_pp1_iter121;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter123_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter123 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter123 <= ap_enable_reg_pp1_iter122;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter124_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter124 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter124 <= ap_enable_reg_pp1_iter123;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter125_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter125 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter125 <= ap_enable_reg_pp1_iter124;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter126_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter126 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter126 <= ap_enable_reg_pp1_iter125;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter127_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter127 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter127 <= ap_enable_reg_pp1_iter126;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter128_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter128 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter128 <= ap_enable_reg_pp1_iter127;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter129_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter129 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter129 <= ap_enable_reg_pp1_iter128;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter13_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter13 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter13 <= ap_enable_reg_pp1_iter12;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter130_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter130 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter130 <= ap_enable_reg_pp1_iter129;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter131_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter131 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter131 <= ap_enable_reg_pp1_iter130;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter132_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter132 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter132 <= ap_enable_reg_pp1_iter131;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter133_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter133 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter133 <= ap_enable_reg_pp1_iter132;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter134_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter134 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter134 <= ap_enable_reg_pp1_iter133;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter135_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter135 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter135 <= ap_enable_reg_pp1_iter134;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter136_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter136 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter136 <= ap_enable_reg_pp1_iter135;
                elsif (((ap_const_lv1_1 = ap_CS_fsm_state139))) then 
                    ap_enable_reg_pp1_iter136 <= ap_const_logic_0;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter14_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter14 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter14 <= ap_enable_reg_pp1_iter13;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter15_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter15 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter15 <= ap_enable_reg_pp1_iter14;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter16_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter16 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter16 <= ap_enable_reg_pp1_iter15;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter17_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter17 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter17 <= ap_enable_reg_pp1_iter16;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter18_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter18 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter18 <= ap_enable_reg_pp1_iter17;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter19_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter19 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter19 <= ap_enable_reg_pp1_iter18;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter2_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter2 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter2 <= ap_enable_reg_pp1_iter1;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter20_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter20 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter20 <= ap_enable_reg_pp1_iter19;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter21_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter21 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter21 <= ap_enable_reg_pp1_iter20;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter22_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter22 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter22 <= ap_enable_reg_pp1_iter21;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter23_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter23 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter23 <= ap_enable_reg_pp1_iter22;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter24_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter24 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter24 <= ap_enable_reg_pp1_iter23;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter25_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter25 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter25 <= ap_enable_reg_pp1_iter24;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter26_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter26 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter26 <= ap_enable_reg_pp1_iter25;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter27_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter27 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter27 <= ap_enable_reg_pp1_iter26;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter28_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter28 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter28 <= ap_enable_reg_pp1_iter27;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter29_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter29 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter29 <= ap_enable_reg_pp1_iter28;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter3_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter3 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter3 <= ap_enable_reg_pp1_iter2;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter30_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter30 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter30 <= ap_enable_reg_pp1_iter29;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter31_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter31 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter31 <= ap_enable_reg_pp1_iter30;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter32_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter32 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter32 <= ap_enable_reg_pp1_iter31;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter33_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter33 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter33 <= ap_enable_reg_pp1_iter32;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter34_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter34 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter34 <= ap_enable_reg_pp1_iter33;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter35_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter35 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter35 <= ap_enable_reg_pp1_iter34;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter36_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter36 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter36 <= ap_enable_reg_pp1_iter35;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter37_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter37 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter37 <= ap_enable_reg_pp1_iter36;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter38_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter38 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter38 <= ap_enable_reg_pp1_iter37;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter39_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter39 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter39 <= ap_enable_reg_pp1_iter38;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter4_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter4 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter4 <= ap_enable_reg_pp1_iter3;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter40_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter40 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter40 <= ap_enable_reg_pp1_iter39;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter41_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter41 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter41 <= ap_enable_reg_pp1_iter40;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter42_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter42 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter42 <= ap_enable_reg_pp1_iter41;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter43_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter43 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter43 <= ap_enable_reg_pp1_iter42;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter44_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter44 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter44 <= ap_enable_reg_pp1_iter43;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter45_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter45 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter45 <= ap_enable_reg_pp1_iter44;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter46_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter46 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter46 <= ap_enable_reg_pp1_iter45;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter47_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter47 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter47 <= ap_enable_reg_pp1_iter46;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter48_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter48 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter48 <= ap_enable_reg_pp1_iter47;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter49_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter49 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter49 <= ap_enable_reg_pp1_iter48;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter5_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter5 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter5 <= ap_enable_reg_pp1_iter4;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter50_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter50 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter50 <= ap_enable_reg_pp1_iter49;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter51_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter51 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter51 <= ap_enable_reg_pp1_iter50;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter52_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter52 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter52 <= ap_enable_reg_pp1_iter51;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter53_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter53 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter53 <= ap_enable_reg_pp1_iter52;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter54_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter54 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter54 <= ap_enable_reg_pp1_iter53;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter55_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter55 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter55 <= ap_enable_reg_pp1_iter54;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter56_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter56 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter56 <= ap_enable_reg_pp1_iter55;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter57_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter57 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter57 <= ap_enable_reg_pp1_iter56;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter58_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter58 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter58 <= ap_enable_reg_pp1_iter57;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter59_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter59 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter59 <= ap_enable_reg_pp1_iter58;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter6_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter6 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter6 <= ap_enable_reg_pp1_iter5;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter60_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter60 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter60 <= ap_enable_reg_pp1_iter59;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter61_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter61 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter61 <= ap_enable_reg_pp1_iter60;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter62_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter62 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter62 <= ap_enable_reg_pp1_iter61;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter63_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter63 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter63 <= ap_enable_reg_pp1_iter62;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter64_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter64 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter64 <= ap_enable_reg_pp1_iter63;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter65_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter65 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter65 <= ap_enable_reg_pp1_iter64;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter66_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter66 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter66 <= ap_enable_reg_pp1_iter65;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter67_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter67 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter67 <= ap_enable_reg_pp1_iter66;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter68_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter68 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter68 <= ap_enable_reg_pp1_iter67;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter69_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter69 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter69 <= ap_enable_reg_pp1_iter68;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter7_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter7 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter7 <= ap_enable_reg_pp1_iter6;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter70_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter70 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter70 <= ap_enable_reg_pp1_iter69;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter71_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter71 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter71 <= ap_enable_reg_pp1_iter70;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter72_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter72 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter72 <= ap_enable_reg_pp1_iter71;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter73_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter73 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter73 <= ap_enable_reg_pp1_iter72;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter74_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter74 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter74 <= ap_enable_reg_pp1_iter73;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter75_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter75 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter75 <= ap_enable_reg_pp1_iter74;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter76_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter76 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter76 <= ap_enable_reg_pp1_iter75;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter77_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter77 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter77 <= ap_enable_reg_pp1_iter76;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter78_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter78 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter78 <= ap_enable_reg_pp1_iter77;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter79_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter79 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter79 <= ap_enable_reg_pp1_iter78;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter8_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter8 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter8 <= ap_enable_reg_pp1_iter7;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter80_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter80 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter80 <= ap_enable_reg_pp1_iter79;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter81_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter81 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter81 <= ap_enable_reg_pp1_iter80;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter82_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter82 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter82 <= ap_enable_reg_pp1_iter81;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter83_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter83 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter83 <= ap_enable_reg_pp1_iter82;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter84_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter84 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter84 <= ap_enable_reg_pp1_iter83;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter85_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter85 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter85 <= ap_enable_reg_pp1_iter84;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter86_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter86 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter86 <= ap_enable_reg_pp1_iter85;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter87_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter87 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter87 <= ap_enable_reg_pp1_iter86;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter88_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter88 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter88 <= ap_enable_reg_pp1_iter87;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter89_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter89 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter89 <= ap_enable_reg_pp1_iter88;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter9_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter9 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter9 <= ap_enable_reg_pp1_iter8;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter90_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter90 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter90 <= ap_enable_reg_pp1_iter89;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter91_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter91 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter91 <= ap_enable_reg_pp1_iter90;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter92_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter92 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter92 <= ap_enable_reg_pp1_iter91;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter93_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter93 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter93 <= ap_enable_reg_pp1_iter92;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter94_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter94 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter94 <= ap_enable_reg_pp1_iter93;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter95_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter95 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter95 <= ap_enable_reg_pp1_iter94;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter96_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter96 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter96 <= ap_enable_reg_pp1_iter95;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter97_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter97 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter97 <= ap_enable_reg_pp1_iter96;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter98_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter98 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter98 <= ap_enable_reg_pp1_iter97;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp1_iter99_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp1_iter99 <= ap_const_logic_0;
            else
                if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then 
                    ap_enable_reg_pp1_iter99 <= ap_enable_reg_pp1_iter98;
                end if; 
            end if;
        end if;
    end process;


    ap_reg_ioackin_gmem_ARREADY_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_reg_ioackin_gmem_ARREADY <= ap_const_logic_0;
            else
                if ((((ap_const_lv1_1 = ap_CS_fsm_pp0_stage0) and (ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) or ((ap_const_lv1_1 = ap_CS_fsm_pp1_stage0) and (ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))))) then 
                    ap_reg_ioackin_gmem_ARREADY <= ap_const_logic_0;
                elsif ((((ap_const_lv1_1 = ap_CS_fsm_pp0_stage0) and (ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_1 = gmem_ARREADY) and not(((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))) or ((ap_const_lv1_1 = ap_CS_fsm_pp1_stage0) and (ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_1 = gmem_ARREADY) and not(((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))))) then 
                    ap_reg_ioackin_gmem_ARREADY <= ap_const_logic_1;
                end if; 
            end if;
        end if;
    end process;


    ap_reg_ioackin_gmem_AWREADY_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_reg_ioackin_gmem_AWREADY <= ap_const_logic_0;
            else
                if ((ap_const_lv1_1 = ap_CS_fsm_state278)) then
                    if (not((ap_const_logic_0 = ap_sig_ioackin_gmem_AWREADY))) then 
                        ap_reg_ioackin_gmem_AWREADY <= ap_const_logic_0;
                    elsif ((ap_const_logic_1 = gmem_AWREADY)) then 
                        ap_reg_ioackin_gmem_AWREADY <= ap_const_logic_1;
                    end if;
                end if; 
            end if;
        end if;
    end process;


    ap_reg_ioackin_gmem_WREADY_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_reg_ioackin_gmem_WREADY <= ap_const_logic_0;
            else
                if ((ap_const_lv1_1 = ap_CS_fsm_state285)) then
                    if (not((ap_const_logic_0 = ap_sig_ioackin_gmem_WREADY))) then 
                        ap_reg_ioackin_gmem_WREADY <= ap_const_logic_0;
                    elsif ((ap_const_logic_1 = gmem_WREADY)) then 
                        ap_reg_ioackin_gmem_WREADY <= ap_const_logic_1;
                    end if;
                end if; 
            end if;
        end if;
    end process;


    indvar7_reg_203_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_lv1_1 = ap_CS_fsm_state139))) then 
                indvar7_reg_203 <= ap_const_lv5_0;
            elsif (((ap_const_lv1_1 = ap_CS_fsm_pp1_stage0) and (ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_lv1_0 = exitcond9_reg_485))) then 
                indvar7_reg_203 <= indvar_next8_reg_489;
            end if; 
        end if;
    end process;

    indvar_reg2mem44_0_i_reg_215_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_lv1_1 = ap_CS_fsm_state278) and not((ap_const_logic_0 = ap_sig_ioackin_gmem_AWREADY)))) then 
                indvar_reg2mem44_0_i_reg_215 <= ap_const_lv5_0;
            elsif (((ap_const_lv1_1 = ap_CS_fsm_state285) and not((ap_const_logic_0 = ap_sig_ioackin_gmem_WREADY)))) then 
                indvar_reg2mem44_0_i_reg_215 <= indvar_inc_reg2mem_reg_511;
            end if; 
        end if;
    end process;

    indvar_reg_191_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_CS_fsm_state1 = ap_const_lv1_1) and not((ap_start = ap_const_logic_0)))) then 
                indvar_reg_191 <= ap_const_lv5_0;
            elsif (((ap_const_lv1_1 = ap_CS_fsm_pp0_stage0) and (ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_lv1_0 = exitcond_reg_472))) then 
                indvar_reg_191 <= indvar_next_reg_476;
            end if; 
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) then
                ap_pipeline_reg_pp0_iter100_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter99_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter100_indvar_reg_191 <= ap_pipeline_reg_pp0_iter99_indvar_reg_191;
                ap_pipeline_reg_pp0_iter101_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter100_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter101_indvar_reg_191 <= ap_pipeline_reg_pp0_iter100_indvar_reg_191;
                ap_pipeline_reg_pp0_iter102_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter101_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter102_indvar_reg_191 <= ap_pipeline_reg_pp0_iter101_indvar_reg_191;
                ap_pipeline_reg_pp0_iter103_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter102_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter103_indvar_reg_191 <= ap_pipeline_reg_pp0_iter102_indvar_reg_191;
                ap_pipeline_reg_pp0_iter104_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter103_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter104_indvar_reg_191 <= ap_pipeline_reg_pp0_iter103_indvar_reg_191;
                ap_pipeline_reg_pp0_iter105_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter104_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter105_indvar_reg_191 <= ap_pipeline_reg_pp0_iter104_indvar_reg_191;
                ap_pipeline_reg_pp0_iter106_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter105_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter106_indvar_reg_191 <= ap_pipeline_reg_pp0_iter105_indvar_reg_191;
                ap_pipeline_reg_pp0_iter107_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter106_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter107_indvar_reg_191 <= ap_pipeline_reg_pp0_iter106_indvar_reg_191;
                ap_pipeline_reg_pp0_iter108_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter107_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter108_indvar_reg_191 <= ap_pipeline_reg_pp0_iter107_indvar_reg_191;
                ap_pipeline_reg_pp0_iter109_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter108_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter109_indvar_reg_191 <= ap_pipeline_reg_pp0_iter108_indvar_reg_191;
                ap_pipeline_reg_pp0_iter10_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter9_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter10_indvar_reg_191 <= ap_pipeline_reg_pp0_iter9_indvar_reg_191;
                ap_pipeline_reg_pp0_iter110_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter109_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter110_indvar_reg_191 <= ap_pipeline_reg_pp0_iter109_indvar_reg_191;
                ap_pipeline_reg_pp0_iter111_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter110_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter111_indvar_reg_191 <= ap_pipeline_reg_pp0_iter110_indvar_reg_191;
                ap_pipeline_reg_pp0_iter112_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter111_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter112_indvar_reg_191 <= ap_pipeline_reg_pp0_iter111_indvar_reg_191;
                ap_pipeline_reg_pp0_iter113_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter112_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter113_indvar_reg_191 <= ap_pipeline_reg_pp0_iter112_indvar_reg_191;
                ap_pipeline_reg_pp0_iter114_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter113_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter114_indvar_reg_191 <= ap_pipeline_reg_pp0_iter113_indvar_reg_191;
                ap_pipeline_reg_pp0_iter115_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter114_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter115_indvar_reg_191 <= ap_pipeline_reg_pp0_iter114_indvar_reg_191;
                ap_pipeline_reg_pp0_iter116_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter115_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter116_indvar_reg_191 <= ap_pipeline_reg_pp0_iter115_indvar_reg_191;
                ap_pipeline_reg_pp0_iter117_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter116_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter117_indvar_reg_191 <= ap_pipeline_reg_pp0_iter116_indvar_reg_191;
                ap_pipeline_reg_pp0_iter118_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter117_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter118_indvar_reg_191 <= ap_pipeline_reg_pp0_iter117_indvar_reg_191;
                ap_pipeline_reg_pp0_iter119_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter118_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter119_indvar_reg_191 <= ap_pipeline_reg_pp0_iter118_indvar_reg_191;
                ap_pipeline_reg_pp0_iter11_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter10_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter11_indvar_reg_191 <= ap_pipeline_reg_pp0_iter10_indvar_reg_191;
                ap_pipeline_reg_pp0_iter120_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter119_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter120_indvar_reg_191 <= ap_pipeline_reg_pp0_iter119_indvar_reg_191;
                ap_pipeline_reg_pp0_iter121_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter120_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter121_indvar_reg_191 <= ap_pipeline_reg_pp0_iter120_indvar_reg_191;
                ap_pipeline_reg_pp0_iter122_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter121_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter122_indvar_reg_191 <= ap_pipeline_reg_pp0_iter121_indvar_reg_191;
                ap_pipeline_reg_pp0_iter123_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter122_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter123_indvar_reg_191 <= ap_pipeline_reg_pp0_iter122_indvar_reg_191;
                ap_pipeline_reg_pp0_iter124_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter123_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter124_indvar_reg_191 <= ap_pipeline_reg_pp0_iter123_indvar_reg_191;
                ap_pipeline_reg_pp0_iter125_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter124_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter125_indvar_reg_191 <= ap_pipeline_reg_pp0_iter124_indvar_reg_191;
                ap_pipeline_reg_pp0_iter126_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter125_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter126_indvar_reg_191 <= ap_pipeline_reg_pp0_iter125_indvar_reg_191;
                ap_pipeline_reg_pp0_iter127_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter126_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter127_indvar_reg_191 <= ap_pipeline_reg_pp0_iter126_indvar_reg_191;
                ap_pipeline_reg_pp0_iter128_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter127_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter128_indvar_reg_191 <= ap_pipeline_reg_pp0_iter127_indvar_reg_191;
                ap_pipeline_reg_pp0_iter129_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter128_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter129_indvar_reg_191 <= ap_pipeline_reg_pp0_iter128_indvar_reg_191;
                ap_pipeline_reg_pp0_iter12_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter11_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter12_indvar_reg_191 <= ap_pipeline_reg_pp0_iter11_indvar_reg_191;
                ap_pipeline_reg_pp0_iter130_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter129_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter130_indvar_reg_191 <= ap_pipeline_reg_pp0_iter129_indvar_reg_191;
                ap_pipeline_reg_pp0_iter131_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter130_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter131_indvar_reg_191 <= ap_pipeline_reg_pp0_iter130_indvar_reg_191;
                ap_pipeline_reg_pp0_iter132_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter131_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter132_indvar_reg_191 <= ap_pipeline_reg_pp0_iter131_indvar_reg_191;
                ap_pipeline_reg_pp0_iter133_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter132_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter133_indvar_reg_191 <= ap_pipeline_reg_pp0_iter132_indvar_reg_191;
                ap_pipeline_reg_pp0_iter134_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter133_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter134_indvar_reg_191 <= ap_pipeline_reg_pp0_iter133_indvar_reg_191;
                ap_pipeline_reg_pp0_iter135_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter134_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter135_indvar_reg_191 <= ap_pipeline_reg_pp0_iter134_indvar_reg_191;
                ap_pipeline_reg_pp0_iter13_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter12_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter13_indvar_reg_191 <= ap_pipeline_reg_pp0_iter12_indvar_reg_191;
                ap_pipeline_reg_pp0_iter14_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter13_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter14_indvar_reg_191 <= ap_pipeline_reg_pp0_iter13_indvar_reg_191;
                ap_pipeline_reg_pp0_iter15_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter14_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter15_indvar_reg_191 <= ap_pipeline_reg_pp0_iter14_indvar_reg_191;
                ap_pipeline_reg_pp0_iter16_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter15_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter16_indvar_reg_191 <= ap_pipeline_reg_pp0_iter15_indvar_reg_191;
                ap_pipeline_reg_pp0_iter17_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter16_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter17_indvar_reg_191 <= ap_pipeline_reg_pp0_iter16_indvar_reg_191;
                ap_pipeline_reg_pp0_iter18_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter17_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter18_indvar_reg_191 <= ap_pipeline_reg_pp0_iter17_indvar_reg_191;
                ap_pipeline_reg_pp0_iter19_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter18_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter19_indvar_reg_191 <= ap_pipeline_reg_pp0_iter18_indvar_reg_191;
                ap_pipeline_reg_pp0_iter20_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter19_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter20_indvar_reg_191 <= ap_pipeline_reg_pp0_iter19_indvar_reg_191;
                ap_pipeline_reg_pp0_iter21_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter20_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter21_indvar_reg_191 <= ap_pipeline_reg_pp0_iter20_indvar_reg_191;
                ap_pipeline_reg_pp0_iter22_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter21_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter22_indvar_reg_191 <= ap_pipeline_reg_pp0_iter21_indvar_reg_191;
                ap_pipeline_reg_pp0_iter23_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter22_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter23_indvar_reg_191 <= ap_pipeline_reg_pp0_iter22_indvar_reg_191;
                ap_pipeline_reg_pp0_iter24_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter23_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter24_indvar_reg_191 <= ap_pipeline_reg_pp0_iter23_indvar_reg_191;
                ap_pipeline_reg_pp0_iter25_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter24_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter25_indvar_reg_191 <= ap_pipeline_reg_pp0_iter24_indvar_reg_191;
                ap_pipeline_reg_pp0_iter26_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter25_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter26_indvar_reg_191 <= ap_pipeline_reg_pp0_iter25_indvar_reg_191;
                ap_pipeline_reg_pp0_iter27_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter26_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter27_indvar_reg_191 <= ap_pipeline_reg_pp0_iter26_indvar_reg_191;
                ap_pipeline_reg_pp0_iter28_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter27_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter28_indvar_reg_191 <= ap_pipeline_reg_pp0_iter27_indvar_reg_191;
                ap_pipeline_reg_pp0_iter29_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter28_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter29_indvar_reg_191 <= ap_pipeline_reg_pp0_iter28_indvar_reg_191;
                ap_pipeline_reg_pp0_iter2_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter1_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter2_indvar_reg_191 <= ap_pipeline_reg_pp0_iter1_indvar_reg_191;
                ap_pipeline_reg_pp0_iter30_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter29_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter30_indvar_reg_191 <= ap_pipeline_reg_pp0_iter29_indvar_reg_191;
                ap_pipeline_reg_pp0_iter31_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter30_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter31_indvar_reg_191 <= ap_pipeline_reg_pp0_iter30_indvar_reg_191;
                ap_pipeline_reg_pp0_iter32_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter31_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter32_indvar_reg_191 <= ap_pipeline_reg_pp0_iter31_indvar_reg_191;
                ap_pipeline_reg_pp0_iter33_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter32_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter33_indvar_reg_191 <= ap_pipeline_reg_pp0_iter32_indvar_reg_191;
                ap_pipeline_reg_pp0_iter34_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter33_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter34_indvar_reg_191 <= ap_pipeline_reg_pp0_iter33_indvar_reg_191;
                ap_pipeline_reg_pp0_iter35_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter34_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter35_indvar_reg_191 <= ap_pipeline_reg_pp0_iter34_indvar_reg_191;
                ap_pipeline_reg_pp0_iter36_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter35_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter36_indvar_reg_191 <= ap_pipeline_reg_pp0_iter35_indvar_reg_191;
                ap_pipeline_reg_pp0_iter37_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter36_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter37_indvar_reg_191 <= ap_pipeline_reg_pp0_iter36_indvar_reg_191;
                ap_pipeline_reg_pp0_iter38_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter37_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter38_indvar_reg_191 <= ap_pipeline_reg_pp0_iter37_indvar_reg_191;
                ap_pipeline_reg_pp0_iter39_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter38_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter39_indvar_reg_191 <= ap_pipeline_reg_pp0_iter38_indvar_reg_191;
                ap_pipeline_reg_pp0_iter3_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter2_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter3_indvar_reg_191 <= ap_pipeline_reg_pp0_iter2_indvar_reg_191;
                ap_pipeline_reg_pp0_iter40_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter39_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter40_indvar_reg_191 <= ap_pipeline_reg_pp0_iter39_indvar_reg_191;
                ap_pipeline_reg_pp0_iter41_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter40_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter41_indvar_reg_191 <= ap_pipeline_reg_pp0_iter40_indvar_reg_191;
                ap_pipeline_reg_pp0_iter42_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter41_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter42_indvar_reg_191 <= ap_pipeline_reg_pp0_iter41_indvar_reg_191;
                ap_pipeline_reg_pp0_iter43_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter42_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter43_indvar_reg_191 <= ap_pipeline_reg_pp0_iter42_indvar_reg_191;
                ap_pipeline_reg_pp0_iter44_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter43_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter44_indvar_reg_191 <= ap_pipeline_reg_pp0_iter43_indvar_reg_191;
                ap_pipeline_reg_pp0_iter45_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter44_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter45_indvar_reg_191 <= ap_pipeline_reg_pp0_iter44_indvar_reg_191;
                ap_pipeline_reg_pp0_iter46_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter45_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter46_indvar_reg_191 <= ap_pipeline_reg_pp0_iter45_indvar_reg_191;
                ap_pipeline_reg_pp0_iter47_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter46_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter47_indvar_reg_191 <= ap_pipeline_reg_pp0_iter46_indvar_reg_191;
                ap_pipeline_reg_pp0_iter48_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter47_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter48_indvar_reg_191 <= ap_pipeline_reg_pp0_iter47_indvar_reg_191;
                ap_pipeline_reg_pp0_iter49_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter48_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter49_indvar_reg_191 <= ap_pipeline_reg_pp0_iter48_indvar_reg_191;
                ap_pipeline_reg_pp0_iter4_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter3_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter4_indvar_reg_191 <= ap_pipeline_reg_pp0_iter3_indvar_reg_191;
                ap_pipeline_reg_pp0_iter50_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter49_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter50_indvar_reg_191 <= ap_pipeline_reg_pp0_iter49_indvar_reg_191;
                ap_pipeline_reg_pp0_iter51_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter50_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter51_indvar_reg_191 <= ap_pipeline_reg_pp0_iter50_indvar_reg_191;
                ap_pipeline_reg_pp0_iter52_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter51_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter52_indvar_reg_191 <= ap_pipeline_reg_pp0_iter51_indvar_reg_191;
                ap_pipeline_reg_pp0_iter53_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter52_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter53_indvar_reg_191 <= ap_pipeline_reg_pp0_iter52_indvar_reg_191;
                ap_pipeline_reg_pp0_iter54_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter53_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter54_indvar_reg_191 <= ap_pipeline_reg_pp0_iter53_indvar_reg_191;
                ap_pipeline_reg_pp0_iter55_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter54_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter55_indvar_reg_191 <= ap_pipeline_reg_pp0_iter54_indvar_reg_191;
                ap_pipeline_reg_pp0_iter56_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter55_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter56_indvar_reg_191 <= ap_pipeline_reg_pp0_iter55_indvar_reg_191;
                ap_pipeline_reg_pp0_iter57_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter56_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter57_indvar_reg_191 <= ap_pipeline_reg_pp0_iter56_indvar_reg_191;
                ap_pipeline_reg_pp0_iter58_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter57_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter58_indvar_reg_191 <= ap_pipeline_reg_pp0_iter57_indvar_reg_191;
                ap_pipeline_reg_pp0_iter59_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter58_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter59_indvar_reg_191 <= ap_pipeline_reg_pp0_iter58_indvar_reg_191;
                ap_pipeline_reg_pp0_iter5_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter4_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter5_indvar_reg_191 <= ap_pipeline_reg_pp0_iter4_indvar_reg_191;
                ap_pipeline_reg_pp0_iter60_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter59_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter60_indvar_reg_191 <= ap_pipeline_reg_pp0_iter59_indvar_reg_191;
                ap_pipeline_reg_pp0_iter61_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter60_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter61_indvar_reg_191 <= ap_pipeline_reg_pp0_iter60_indvar_reg_191;
                ap_pipeline_reg_pp0_iter62_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter61_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter62_indvar_reg_191 <= ap_pipeline_reg_pp0_iter61_indvar_reg_191;
                ap_pipeline_reg_pp0_iter63_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter62_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter63_indvar_reg_191 <= ap_pipeline_reg_pp0_iter62_indvar_reg_191;
                ap_pipeline_reg_pp0_iter64_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter63_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter64_indvar_reg_191 <= ap_pipeline_reg_pp0_iter63_indvar_reg_191;
                ap_pipeline_reg_pp0_iter65_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter64_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter65_indvar_reg_191 <= ap_pipeline_reg_pp0_iter64_indvar_reg_191;
                ap_pipeline_reg_pp0_iter66_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter65_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter66_indvar_reg_191 <= ap_pipeline_reg_pp0_iter65_indvar_reg_191;
                ap_pipeline_reg_pp0_iter67_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter66_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter67_indvar_reg_191 <= ap_pipeline_reg_pp0_iter66_indvar_reg_191;
                ap_pipeline_reg_pp0_iter68_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter67_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter68_indvar_reg_191 <= ap_pipeline_reg_pp0_iter67_indvar_reg_191;
                ap_pipeline_reg_pp0_iter69_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter68_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter69_indvar_reg_191 <= ap_pipeline_reg_pp0_iter68_indvar_reg_191;
                ap_pipeline_reg_pp0_iter6_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter5_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter6_indvar_reg_191 <= ap_pipeline_reg_pp0_iter5_indvar_reg_191;
                ap_pipeline_reg_pp0_iter70_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter69_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter70_indvar_reg_191 <= ap_pipeline_reg_pp0_iter69_indvar_reg_191;
                ap_pipeline_reg_pp0_iter71_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter70_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter71_indvar_reg_191 <= ap_pipeline_reg_pp0_iter70_indvar_reg_191;
                ap_pipeline_reg_pp0_iter72_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter71_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter72_indvar_reg_191 <= ap_pipeline_reg_pp0_iter71_indvar_reg_191;
                ap_pipeline_reg_pp0_iter73_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter72_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter73_indvar_reg_191 <= ap_pipeline_reg_pp0_iter72_indvar_reg_191;
                ap_pipeline_reg_pp0_iter74_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter73_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter74_indvar_reg_191 <= ap_pipeline_reg_pp0_iter73_indvar_reg_191;
                ap_pipeline_reg_pp0_iter75_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter74_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter75_indvar_reg_191 <= ap_pipeline_reg_pp0_iter74_indvar_reg_191;
                ap_pipeline_reg_pp0_iter76_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter75_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter76_indvar_reg_191 <= ap_pipeline_reg_pp0_iter75_indvar_reg_191;
                ap_pipeline_reg_pp0_iter77_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter76_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter77_indvar_reg_191 <= ap_pipeline_reg_pp0_iter76_indvar_reg_191;
                ap_pipeline_reg_pp0_iter78_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter77_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter78_indvar_reg_191 <= ap_pipeline_reg_pp0_iter77_indvar_reg_191;
                ap_pipeline_reg_pp0_iter79_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter78_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter79_indvar_reg_191 <= ap_pipeline_reg_pp0_iter78_indvar_reg_191;
                ap_pipeline_reg_pp0_iter7_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter6_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter7_indvar_reg_191 <= ap_pipeline_reg_pp0_iter6_indvar_reg_191;
                ap_pipeline_reg_pp0_iter80_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter79_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter80_indvar_reg_191 <= ap_pipeline_reg_pp0_iter79_indvar_reg_191;
                ap_pipeline_reg_pp0_iter81_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter80_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter81_indvar_reg_191 <= ap_pipeline_reg_pp0_iter80_indvar_reg_191;
                ap_pipeline_reg_pp0_iter82_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter81_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter82_indvar_reg_191 <= ap_pipeline_reg_pp0_iter81_indvar_reg_191;
                ap_pipeline_reg_pp0_iter83_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter82_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter83_indvar_reg_191 <= ap_pipeline_reg_pp0_iter82_indvar_reg_191;
                ap_pipeline_reg_pp0_iter84_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter83_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter84_indvar_reg_191 <= ap_pipeline_reg_pp0_iter83_indvar_reg_191;
                ap_pipeline_reg_pp0_iter85_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter84_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter85_indvar_reg_191 <= ap_pipeline_reg_pp0_iter84_indvar_reg_191;
                ap_pipeline_reg_pp0_iter86_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter85_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter86_indvar_reg_191 <= ap_pipeline_reg_pp0_iter85_indvar_reg_191;
                ap_pipeline_reg_pp0_iter87_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter86_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter87_indvar_reg_191 <= ap_pipeline_reg_pp0_iter86_indvar_reg_191;
                ap_pipeline_reg_pp0_iter88_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter87_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter88_indvar_reg_191 <= ap_pipeline_reg_pp0_iter87_indvar_reg_191;
                ap_pipeline_reg_pp0_iter89_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter88_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter89_indvar_reg_191 <= ap_pipeline_reg_pp0_iter88_indvar_reg_191;
                ap_pipeline_reg_pp0_iter8_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter7_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter8_indvar_reg_191 <= ap_pipeline_reg_pp0_iter7_indvar_reg_191;
                ap_pipeline_reg_pp0_iter90_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter89_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter90_indvar_reg_191 <= ap_pipeline_reg_pp0_iter89_indvar_reg_191;
                ap_pipeline_reg_pp0_iter91_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter90_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter91_indvar_reg_191 <= ap_pipeline_reg_pp0_iter90_indvar_reg_191;
                ap_pipeline_reg_pp0_iter92_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter91_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter92_indvar_reg_191 <= ap_pipeline_reg_pp0_iter91_indvar_reg_191;
                ap_pipeline_reg_pp0_iter93_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter92_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter93_indvar_reg_191 <= ap_pipeline_reg_pp0_iter92_indvar_reg_191;
                ap_pipeline_reg_pp0_iter94_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter93_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter94_indvar_reg_191 <= ap_pipeline_reg_pp0_iter93_indvar_reg_191;
                ap_pipeline_reg_pp0_iter95_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter94_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter95_indvar_reg_191 <= ap_pipeline_reg_pp0_iter94_indvar_reg_191;
                ap_pipeline_reg_pp0_iter96_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter95_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter96_indvar_reg_191 <= ap_pipeline_reg_pp0_iter95_indvar_reg_191;
                ap_pipeline_reg_pp0_iter97_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter96_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter97_indvar_reg_191 <= ap_pipeline_reg_pp0_iter96_indvar_reg_191;
                ap_pipeline_reg_pp0_iter98_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter97_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter98_indvar_reg_191 <= ap_pipeline_reg_pp0_iter97_indvar_reg_191;
                ap_pipeline_reg_pp0_iter99_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter98_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter99_indvar_reg_191 <= ap_pipeline_reg_pp0_iter98_indvar_reg_191;
                ap_pipeline_reg_pp0_iter9_exitcond_reg_472 <= ap_pipeline_reg_pp0_iter8_exitcond_reg_472;
                ap_pipeline_reg_pp0_iter9_indvar_reg_191 <= ap_pipeline_reg_pp0_iter8_indvar_reg_191;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_lv1_1 = ap_CS_fsm_pp0_stage0) and not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))))) then
                ap_pipeline_reg_pp0_iter1_exitcond_reg_472 <= exitcond_reg_472;
                ap_pipeline_reg_pp0_iter1_indvar_reg_191 <= indvar_reg_191;
                exitcond_reg_472 <= exitcond_fu_308_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))) then
                ap_pipeline_reg_pp1_iter100_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter99_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter100_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter99_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter101_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter100_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter101_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter100_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter102_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter101_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter102_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter101_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter103_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter102_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter103_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter102_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter104_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter103_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter104_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter103_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter105_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter104_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter105_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter104_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter106_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter105_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter106_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter105_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter107_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter106_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter107_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter106_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter108_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter107_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter108_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter107_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter109_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter108_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter109_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter108_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter10_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter9_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter10_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter9_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter110_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter109_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter110_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter109_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter111_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter110_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter111_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter110_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter112_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter111_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter112_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter111_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter113_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter112_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter113_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter112_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter114_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter113_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter114_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter113_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter115_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter114_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter115_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter114_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter116_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter115_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter116_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter115_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter117_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter116_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter117_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter116_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter118_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter117_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter118_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter117_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter119_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter118_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter119_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter118_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter11_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter10_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter11_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter10_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter120_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter119_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter120_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter119_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter121_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter120_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter121_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter120_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter122_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter121_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter122_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter121_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter123_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter122_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter123_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter122_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter124_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter123_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter124_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter123_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter125_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter124_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter125_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter124_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter126_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter125_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter126_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter125_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter127_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter126_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter127_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter126_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter128_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter127_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter128_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter127_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter129_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter128_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter129_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter128_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter12_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter11_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter12_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter11_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter130_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter129_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter130_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter129_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter131_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter130_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter131_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter130_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter132_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter131_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter132_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter131_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter133_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter132_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter133_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter132_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter134_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter133_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter134_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter133_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter135_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter134_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter135_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter134_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter13_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter12_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter13_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter12_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter14_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter13_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter14_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter13_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter15_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter14_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter15_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter14_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter16_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter15_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter16_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter15_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter17_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter16_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter17_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter16_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter18_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter17_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter18_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter17_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter19_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter18_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter19_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter18_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter20_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter19_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter20_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter19_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter21_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter20_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter21_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter20_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter22_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter21_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter22_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter21_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter23_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter22_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter23_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter22_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter24_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter23_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter24_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter23_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter25_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter24_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter25_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter24_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter26_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter25_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter26_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter25_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter27_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter26_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter27_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter26_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter28_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter27_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter28_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter27_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter29_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter28_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter29_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter28_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter2_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter1_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter2_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter1_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter30_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter29_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter30_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter29_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter31_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter30_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter31_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter30_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter32_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter31_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter32_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter31_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter33_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter32_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter33_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter32_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter34_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter33_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter34_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter33_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter35_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter34_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter35_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter34_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter36_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter35_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter36_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter35_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter37_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter36_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter37_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter36_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter38_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter37_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter38_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter37_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter39_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter38_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter39_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter38_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter3_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter2_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter3_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter2_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter40_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter39_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter40_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter39_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter41_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter40_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter41_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter40_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter42_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter41_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter42_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter41_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter43_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter42_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter43_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter42_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter44_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter43_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter44_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter43_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter45_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter44_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter45_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter44_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter46_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter45_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter46_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter45_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter47_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter46_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter47_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter46_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter48_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter47_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter48_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter47_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter49_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter48_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter49_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter48_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter4_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter3_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter4_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter3_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter50_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter49_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter50_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter49_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter51_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter50_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter51_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter50_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter52_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter51_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter52_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter51_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter53_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter52_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter53_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter52_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter54_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter53_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter54_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter53_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter55_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter54_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter55_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter54_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter56_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter55_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter56_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter55_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter57_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter56_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter57_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter56_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter58_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter57_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter58_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter57_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter59_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter58_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter59_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter58_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter5_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter4_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter5_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter4_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter60_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter59_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter60_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter59_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter61_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter60_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter61_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter60_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter62_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter61_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter62_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter61_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter63_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter62_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter63_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter62_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter64_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter63_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter64_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter63_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter65_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter64_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter65_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter64_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter66_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter65_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter66_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter65_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter67_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter66_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter67_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter66_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter68_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter67_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter68_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter67_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter69_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter68_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter69_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter68_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter6_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter5_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter6_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter5_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter70_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter69_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter70_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter69_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter71_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter70_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter71_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter70_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter72_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter71_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter72_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter71_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter73_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter72_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter73_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter72_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter74_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter73_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter74_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter73_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter75_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter74_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter75_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter74_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter76_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter75_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter76_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter75_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter77_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter76_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter77_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter76_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter78_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter77_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter78_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter77_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter79_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter78_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter79_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter78_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter7_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter6_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter7_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter6_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter80_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter79_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter80_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter79_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter81_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter80_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter81_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter80_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter82_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter81_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter82_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter81_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter83_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter82_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter83_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter82_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter84_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter83_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter84_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter83_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter85_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter84_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter85_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter84_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter86_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter85_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter86_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter85_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter87_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter86_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter87_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter86_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter88_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter87_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter88_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter87_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter89_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter88_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter89_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter88_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter8_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter7_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter8_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter7_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter90_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter89_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter90_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter89_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter91_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter90_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter91_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter90_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter92_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter91_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter92_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter91_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter93_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter92_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter93_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter92_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter94_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter93_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter94_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter93_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter95_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter94_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter95_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter94_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter96_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter95_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter96_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter95_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter97_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter96_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter97_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter96_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter98_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter97_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter98_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter97_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter99_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter98_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter99_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter98_indvar7_reg_203;
                ap_pipeline_reg_pp1_iter9_exitcond9_reg_485 <= ap_pipeline_reg_pp1_iter8_exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter9_indvar7_reg_203 <= ap_pipeline_reg_pp1_iter8_indvar7_reg_203;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_lv1_1 = ap_CS_fsm_pp1_stage0) and not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))))) then
                ap_pipeline_reg_pp1_iter1_exitcond9_reg_485 <= exitcond9_reg_485;
                ap_pipeline_reg_pp1_iter1_indvar7_reg_203 <= indvar7_reg_203;
                exitcond9_reg_485 <= exitcond9_fu_336_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_CS_fsm_state1 = ap_const_lv1_1) and not((ap_start = ap_const_logic_0)))) then
                    arg_x_reg_455(29 downto 0) <= tmp_10_fu_264_p1(29 downto 0);
                    arg_y_reg_461(29 downto 0) <= tmp_11_fu_284_p1(29 downto 0);
                global_offset_x_read_reg_435 <= global_offset_x;
                tmp_1_reg_445 <= tmp_1_fu_238_p1;
                    tmp_6_cast_reg_467(29 downto 0) <= tmp_6_cast_fu_304_p1(29 downto 0);
                    tmp_cast_reg_450(5 downto 4) <= tmp_cast_fu_246_p3(5 downto 4);
                tmp_reg_440 <= tmp_fu_234_p1;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_lv1_1 = ap_CS_fsm_state279))) then
                indvar_inc_reg2mem_reg_511 <= indvar_inc_reg2mem_fu_405_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_lv1_1 = ap_CS_fsm_pp1_stage0) and not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp1_iter0))) then
                indvar_next8_reg_489 <= indvar_next8_fu_342_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_lv1_1 = ap_CS_fsm_pp0_stage0) and not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp0_iter0))) then
                indvar_next_reg_476 <= indvar_next_fu_314_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_lv1_1 = ap_CS_fsm_pp0_stage0) and not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_lv1_0 = exitcond_fu_308_p2))) then
                isIter0_reg_481 <= isIter0_fu_320_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_lv1_1 = ap_CS_fsm_pp1_stage0) and not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_lv1_0 = exitcond9_fu_336_p2))) then
                isIter_reg_494 <= isIter_fu_348_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))))) then
                reg_230 <= gmem_RDATA;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_lv1_1 = ap_CS_fsm_state277))) then
                tmp_16_reg_498 <= tmp_16_fu_384_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_lv1_1 = ap_CS_fsm_state284))) then
                tmp_3_reg_536 <= grp_fu_226_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_lv1_1 = ap_CS_fsm_state280))) then
                x0_load_reg_526 <= x0_q0;
                y0_load_reg_531 <= y0_q0;
            end if;
        end if;
    end process;
    tmp_cast_reg_450(3 downto 0) <= "0000";
    arg_x_reg_455(31 downto 30) <= "00";
    arg_y_reg_461(31 downto 30) <= "00";
    tmp_6_cast_reg_467(30) <= '0';

    ap_NS_fsm_assign_proc : process (ap_start, ap_CS_fsm, ap_enable_reg_pp0_iter1, isIter0_reg_481, ap_enable_reg_pp0_iter135, ap_pipeline_reg_pp0_iter134_exitcond_reg_472, ap_enable_reg_pp1_iter1, isIter_reg_494, ap_enable_reg_pp1_iter135, ap_pipeline_reg_pp1_iter134_exitcond9_reg_485, gmem_RVALID, gmem_BVALID, ap_sig_ioackin_gmem_ARREADY, exitcond_fu_308_p2, ap_enable_reg_pp0_iter0, exitcond9_fu_336_p2, ap_enable_reg_pp1_iter0, ap_sig_ioackin_gmem_AWREADY, tmp_9_fu_399_p2, ap_enable_reg_pp0_iter136, ap_enable_reg_pp1_iter136, ap_sig_ioackin_gmem_WREADY)
    begin
        case ap_CS_fsm is
            when ap_ST_fsm_state1 => 
                if (not((ap_start = ap_const_logic_0))) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage0;
                else
                    ap_NS_fsm <= ap_ST_fsm_state1;
                end if;
            when ap_ST_fsm_pp0_stage0 => 
                if ((not((not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp0_iter136) and not((ap_const_logic_1 = ap_enable_reg_pp0_iter135)))) and not((not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp0_iter0) and not((ap_const_lv1_0 = exitcond_fu_308_p2)) and not((ap_const_logic_1 = ap_enable_reg_pp0_iter1)))))) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage0;
                elsif (((not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp0_iter136) and not((ap_const_logic_1 = ap_enable_reg_pp0_iter135))) or (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp0_iter0) and not((ap_const_lv1_0 = exitcond_fu_308_p2)) and not((ap_const_logic_1 = ap_enable_reg_pp0_iter1))))) then
                    ap_NS_fsm <= ap_ST_fsm_state139;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage0;
                end if;
            when ap_ST_fsm_state139 => 
                ap_NS_fsm <= ap_ST_fsm_pp1_stage0;
            when ap_ST_fsm_pp1_stage0 => 
                if ((not((not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp1_iter136) and not((ap_const_logic_1 = ap_enable_reg_pp1_iter135)))) and not((not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp1_iter0) and not((ap_const_lv1_0 = exitcond9_fu_336_p2)) and not((ap_const_logic_1 = ap_enable_reg_pp1_iter1)))))) then
                    ap_NS_fsm <= ap_ST_fsm_pp1_stage0;
                elsif (((not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp1_iter136) and not((ap_const_logic_1 = ap_enable_reg_pp1_iter135))) or (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp1_iter0) and not((ap_const_lv1_0 = exitcond9_fu_336_p2)) and not((ap_const_logic_1 = ap_enable_reg_pp1_iter1))))) then
                    ap_NS_fsm <= ap_ST_fsm_state277;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp1_stage0;
                end if;
            when ap_ST_fsm_state277 => 
                ap_NS_fsm <= ap_ST_fsm_state278;
            when ap_ST_fsm_state278 => 
                if (not((ap_const_logic_0 = ap_sig_ioackin_gmem_AWREADY))) then
                    ap_NS_fsm <= ap_ST_fsm_state279;
                else
                    ap_NS_fsm <= ap_ST_fsm_state278;
                end if;
            when ap_ST_fsm_state279 => 
                if (not((ap_const_lv1_0 = tmp_9_fu_399_p2))) then
                    ap_NS_fsm <= ap_ST_fsm_state286;
                else
                    ap_NS_fsm <= ap_ST_fsm_state280;
                end if;
            when ap_ST_fsm_state280 => 
                ap_NS_fsm <= ap_ST_fsm_state281;
            when ap_ST_fsm_state281 => 
                ap_NS_fsm <= ap_ST_fsm_state282;
            when ap_ST_fsm_state282 => 
                ap_NS_fsm <= ap_ST_fsm_state283;
            when ap_ST_fsm_state283 => 
                ap_NS_fsm <= ap_ST_fsm_state284;
            when ap_ST_fsm_state284 => 
                ap_NS_fsm <= ap_ST_fsm_state285;
            when ap_ST_fsm_state285 => 
                if (not((ap_const_logic_0 = ap_sig_ioackin_gmem_WREADY))) then
                    ap_NS_fsm <= ap_ST_fsm_state279;
                else
                    ap_NS_fsm <= ap_ST_fsm_state285;
                end if;
            when ap_ST_fsm_state286 => 
                ap_NS_fsm <= ap_ST_fsm_state287;
            when ap_ST_fsm_state287 => 
                ap_NS_fsm <= ap_ST_fsm_state288;
            when ap_ST_fsm_state288 => 
                ap_NS_fsm <= ap_ST_fsm_state289;
            when ap_ST_fsm_state289 => 
                ap_NS_fsm <= ap_ST_fsm_state290;
            when ap_ST_fsm_state290 => 
                ap_NS_fsm <= ap_ST_fsm_state291;
            when ap_ST_fsm_state291 => 
                ap_NS_fsm <= ap_ST_fsm_state292;
            when ap_ST_fsm_state292 => 
                ap_NS_fsm <= ap_ST_fsm_state293;
            when ap_ST_fsm_state293 => 
                ap_NS_fsm <= ap_ST_fsm_state294;
            when ap_ST_fsm_state294 => 
                ap_NS_fsm <= ap_ST_fsm_state295;
            when ap_ST_fsm_state295 => 
                ap_NS_fsm <= ap_ST_fsm_state296;
            when ap_ST_fsm_state296 => 
                ap_NS_fsm <= ap_ST_fsm_state297;
            when ap_ST_fsm_state297 => 
                ap_NS_fsm <= ap_ST_fsm_state298;
            when ap_ST_fsm_state298 => 
                ap_NS_fsm <= ap_ST_fsm_state299;
            when ap_ST_fsm_state299 => 
                ap_NS_fsm <= ap_ST_fsm_state300;
            when ap_ST_fsm_state300 => 
                ap_NS_fsm <= ap_ST_fsm_state301;
            when ap_ST_fsm_state301 => 
                ap_NS_fsm <= ap_ST_fsm_state302;
            when ap_ST_fsm_state302 => 
                ap_NS_fsm <= ap_ST_fsm_state303;
            when ap_ST_fsm_state303 => 
                ap_NS_fsm <= ap_ST_fsm_state304;
            when ap_ST_fsm_state304 => 
                ap_NS_fsm <= ap_ST_fsm_state305;
            when ap_ST_fsm_state305 => 
                ap_NS_fsm <= ap_ST_fsm_state306;
            when ap_ST_fsm_state306 => 
                ap_NS_fsm <= ap_ST_fsm_state307;
            when ap_ST_fsm_state307 => 
                ap_NS_fsm <= ap_ST_fsm_state308;
            when ap_ST_fsm_state308 => 
                ap_NS_fsm <= ap_ST_fsm_state309;
            when ap_ST_fsm_state309 => 
                ap_NS_fsm <= ap_ST_fsm_state310;
            when ap_ST_fsm_state310 => 
                ap_NS_fsm <= ap_ST_fsm_state311;
            when ap_ST_fsm_state311 => 
                ap_NS_fsm <= ap_ST_fsm_state312;
            when ap_ST_fsm_state312 => 
                ap_NS_fsm <= ap_ST_fsm_state313;
            when ap_ST_fsm_state313 => 
                ap_NS_fsm <= ap_ST_fsm_state314;
            when ap_ST_fsm_state314 => 
                ap_NS_fsm <= ap_ST_fsm_state315;
            when ap_ST_fsm_state315 => 
                ap_NS_fsm <= ap_ST_fsm_state316;
            when ap_ST_fsm_state316 => 
                ap_NS_fsm <= ap_ST_fsm_state317;
            when ap_ST_fsm_state317 => 
                ap_NS_fsm <= ap_ST_fsm_state318;
            when ap_ST_fsm_state318 => 
                ap_NS_fsm <= ap_ST_fsm_state319;
            when ap_ST_fsm_state319 => 
                ap_NS_fsm <= ap_ST_fsm_state320;
            when ap_ST_fsm_state320 => 
                ap_NS_fsm <= ap_ST_fsm_state321;
            when ap_ST_fsm_state321 => 
                ap_NS_fsm <= ap_ST_fsm_state322;
            when ap_ST_fsm_state322 => 
                ap_NS_fsm <= ap_ST_fsm_state323;
            when ap_ST_fsm_state323 => 
                ap_NS_fsm <= ap_ST_fsm_state324;
            when ap_ST_fsm_state324 => 
                ap_NS_fsm <= ap_ST_fsm_state325;
            when ap_ST_fsm_state325 => 
                ap_NS_fsm <= ap_ST_fsm_state326;
            when ap_ST_fsm_state326 => 
                ap_NS_fsm <= ap_ST_fsm_state327;
            when ap_ST_fsm_state327 => 
                ap_NS_fsm <= ap_ST_fsm_state328;
            when ap_ST_fsm_state328 => 
                ap_NS_fsm <= ap_ST_fsm_state329;
            when ap_ST_fsm_state329 => 
                ap_NS_fsm <= ap_ST_fsm_state330;
            when ap_ST_fsm_state330 => 
                ap_NS_fsm <= ap_ST_fsm_state331;
            when ap_ST_fsm_state331 => 
                ap_NS_fsm <= ap_ST_fsm_state332;
            when ap_ST_fsm_state332 => 
                ap_NS_fsm <= ap_ST_fsm_state333;
            when ap_ST_fsm_state333 => 
                ap_NS_fsm <= ap_ST_fsm_state334;
            when ap_ST_fsm_state334 => 
                ap_NS_fsm <= ap_ST_fsm_state335;
            when ap_ST_fsm_state335 => 
                ap_NS_fsm <= ap_ST_fsm_state336;
            when ap_ST_fsm_state336 => 
                ap_NS_fsm <= ap_ST_fsm_state337;
            when ap_ST_fsm_state337 => 
                ap_NS_fsm <= ap_ST_fsm_state338;
            when ap_ST_fsm_state338 => 
                ap_NS_fsm <= ap_ST_fsm_state339;
            when ap_ST_fsm_state339 => 
                ap_NS_fsm <= ap_ST_fsm_state340;
            when ap_ST_fsm_state340 => 
                ap_NS_fsm <= ap_ST_fsm_state341;
            when ap_ST_fsm_state341 => 
                ap_NS_fsm <= ap_ST_fsm_state342;
            when ap_ST_fsm_state342 => 
                ap_NS_fsm <= ap_ST_fsm_state343;
            when ap_ST_fsm_state343 => 
                ap_NS_fsm <= ap_ST_fsm_state344;
            when ap_ST_fsm_state344 => 
                ap_NS_fsm <= ap_ST_fsm_state345;
            when ap_ST_fsm_state345 => 
                ap_NS_fsm <= ap_ST_fsm_state346;
            when ap_ST_fsm_state346 => 
                ap_NS_fsm <= ap_ST_fsm_state347;
            when ap_ST_fsm_state347 => 
                ap_NS_fsm <= ap_ST_fsm_state348;
            when ap_ST_fsm_state348 => 
                ap_NS_fsm <= ap_ST_fsm_state349;
            when ap_ST_fsm_state349 => 
                ap_NS_fsm <= ap_ST_fsm_state350;
            when ap_ST_fsm_state350 => 
                ap_NS_fsm <= ap_ST_fsm_state351;
            when ap_ST_fsm_state351 => 
                ap_NS_fsm <= ap_ST_fsm_state352;
            when ap_ST_fsm_state352 => 
                ap_NS_fsm <= ap_ST_fsm_state353;
            when ap_ST_fsm_state353 => 
                ap_NS_fsm <= ap_ST_fsm_state354;
            when ap_ST_fsm_state354 => 
                ap_NS_fsm <= ap_ST_fsm_state355;
            when ap_ST_fsm_state355 => 
                ap_NS_fsm <= ap_ST_fsm_state356;
            when ap_ST_fsm_state356 => 
                ap_NS_fsm <= ap_ST_fsm_state357;
            when ap_ST_fsm_state357 => 
                ap_NS_fsm <= ap_ST_fsm_state358;
            when ap_ST_fsm_state358 => 
                ap_NS_fsm <= ap_ST_fsm_state359;
            when ap_ST_fsm_state359 => 
                ap_NS_fsm <= ap_ST_fsm_state360;
            when ap_ST_fsm_state360 => 
                ap_NS_fsm <= ap_ST_fsm_state361;
            when ap_ST_fsm_state361 => 
                ap_NS_fsm <= ap_ST_fsm_state362;
            when ap_ST_fsm_state362 => 
                ap_NS_fsm <= ap_ST_fsm_state363;
            when ap_ST_fsm_state363 => 
                ap_NS_fsm <= ap_ST_fsm_state364;
            when ap_ST_fsm_state364 => 
                ap_NS_fsm <= ap_ST_fsm_state365;
            when ap_ST_fsm_state365 => 
                ap_NS_fsm <= ap_ST_fsm_state366;
            when ap_ST_fsm_state366 => 
                ap_NS_fsm <= ap_ST_fsm_state367;
            when ap_ST_fsm_state367 => 
                ap_NS_fsm <= ap_ST_fsm_state368;
            when ap_ST_fsm_state368 => 
                ap_NS_fsm <= ap_ST_fsm_state369;
            when ap_ST_fsm_state369 => 
                ap_NS_fsm <= ap_ST_fsm_state370;
            when ap_ST_fsm_state370 => 
                ap_NS_fsm <= ap_ST_fsm_state371;
            when ap_ST_fsm_state371 => 
                ap_NS_fsm <= ap_ST_fsm_state372;
            when ap_ST_fsm_state372 => 
                ap_NS_fsm <= ap_ST_fsm_state373;
            when ap_ST_fsm_state373 => 
                ap_NS_fsm <= ap_ST_fsm_state374;
            when ap_ST_fsm_state374 => 
                ap_NS_fsm <= ap_ST_fsm_state375;
            when ap_ST_fsm_state375 => 
                ap_NS_fsm <= ap_ST_fsm_state376;
            when ap_ST_fsm_state376 => 
                ap_NS_fsm <= ap_ST_fsm_state377;
            when ap_ST_fsm_state377 => 
                ap_NS_fsm <= ap_ST_fsm_state378;
            when ap_ST_fsm_state378 => 
                ap_NS_fsm <= ap_ST_fsm_state379;
            when ap_ST_fsm_state379 => 
                ap_NS_fsm <= ap_ST_fsm_state380;
            when ap_ST_fsm_state380 => 
                ap_NS_fsm <= ap_ST_fsm_state381;
            when ap_ST_fsm_state381 => 
                ap_NS_fsm <= ap_ST_fsm_state382;
            when ap_ST_fsm_state382 => 
                ap_NS_fsm <= ap_ST_fsm_state383;
            when ap_ST_fsm_state383 => 
                ap_NS_fsm <= ap_ST_fsm_state384;
            when ap_ST_fsm_state384 => 
                ap_NS_fsm <= ap_ST_fsm_state385;
            when ap_ST_fsm_state385 => 
                ap_NS_fsm <= ap_ST_fsm_state386;
            when ap_ST_fsm_state386 => 
                ap_NS_fsm <= ap_ST_fsm_state387;
            when ap_ST_fsm_state387 => 
                ap_NS_fsm <= ap_ST_fsm_state388;
            when ap_ST_fsm_state388 => 
                ap_NS_fsm <= ap_ST_fsm_state389;
            when ap_ST_fsm_state389 => 
                ap_NS_fsm <= ap_ST_fsm_state390;
            when ap_ST_fsm_state390 => 
                ap_NS_fsm <= ap_ST_fsm_state391;
            when ap_ST_fsm_state391 => 
                ap_NS_fsm <= ap_ST_fsm_state392;
            when ap_ST_fsm_state392 => 
                ap_NS_fsm <= ap_ST_fsm_state393;
            when ap_ST_fsm_state393 => 
                ap_NS_fsm <= ap_ST_fsm_state394;
            when ap_ST_fsm_state394 => 
                ap_NS_fsm <= ap_ST_fsm_state395;
            when ap_ST_fsm_state395 => 
                ap_NS_fsm <= ap_ST_fsm_state396;
            when ap_ST_fsm_state396 => 
                ap_NS_fsm <= ap_ST_fsm_state397;
            when ap_ST_fsm_state397 => 
                ap_NS_fsm <= ap_ST_fsm_state398;
            when ap_ST_fsm_state398 => 
                ap_NS_fsm <= ap_ST_fsm_state399;
            when ap_ST_fsm_state399 => 
                ap_NS_fsm <= ap_ST_fsm_state400;
            when ap_ST_fsm_state400 => 
                ap_NS_fsm <= ap_ST_fsm_state401;
            when ap_ST_fsm_state401 => 
                ap_NS_fsm <= ap_ST_fsm_state402;
            when ap_ST_fsm_state402 => 
                ap_NS_fsm <= ap_ST_fsm_state403;
            when ap_ST_fsm_state403 => 
                ap_NS_fsm <= ap_ST_fsm_state404;
            when ap_ST_fsm_state404 => 
                ap_NS_fsm <= ap_ST_fsm_state405;
            when ap_ST_fsm_state405 => 
                ap_NS_fsm <= ap_ST_fsm_state406;
            when ap_ST_fsm_state406 => 
                ap_NS_fsm <= ap_ST_fsm_state407;
            when ap_ST_fsm_state407 => 
                ap_NS_fsm <= ap_ST_fsm_state408;
            when ap_ST_fsm_state408 => 
                ap_NS_fsm <= ap_ST_fsm_state409;
            when ap_ST_fsm_state409 => 
                ap_NS_fsm <= ap_ST_fsm_state410;
            when ap_ST_fsm_state410 => 
                ap_NS_fsm <= ap_ST_fsm_state411;
            when ap_ST_fsm_state411 => 
                ap_NS_fsm <= ap_ST_fsm_state412;
            when ap_ST_fsm_state412 => 
                ap_NS_fsm <= ap_ST_fsm_state413;
            when ap_ST_fsm_state413 => 
                ap_NS_fsm <= ap_ST_fsm_state414;
            when ap_ST_fsm_state414 => 
                ap_NS_fsm <= ap_ST_fsm_state415;
            when ap_ST_fsm_state415 => 
                ap_NS_fsm <= ap_ST_fsm_state416;
            when ap_ST_fsm_state416 => 
                if (not((gmem_BVALID = ap_const_logic_0))) then
                    ap_NS_fsm <= ap_ST_fsm_state1;
                else
                    ap_NS_fsm <= ap_ST_fsm_state416;
                end if;
            when others =>  
                ap_NS_fsm <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
        end case;
    end process;
    ap_CS_fsm_pp0_stage0 <= ap_CS_fsm(1 downto 1);
    ap_CS_fsm_pp1_stage0 <= ap_CS_fsm(3 downto 3);
    ap_CS_fsm_state1 <= ap_CS_fsm(0 downto 0);
    ap_CS_fsm_state139 <= ap_CS_fsm(2 downto 2);
    ap_CS_fsm_state277 <= ap_CS_fsm(4 downto 4);
    ap_CS_fsm_state278 <= ap_CS_fsm(5 downto 5);
    ap_CS_fsm_state279 <= ap_CS_fsm(6 downto 6);
    ap_CS_fsm_state280 <= ap_CS_fsm(7 downto 7);
    ap_CS_fsm_state281 <= ap_CS_fsm(8 downto 8);
    ap_CS_fsm_state284 <= ap_CS_fsm(11 downto 11);
    ap_CS_fsm_state285 <= ap_CS_fsm(12 downto 12);
    ap_CS_fsm_state416 <= ap_CS_fsm(143 downto 143);

    ap_condition_1658_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_enable_reg_pp0_iter1, isIter0_reg_481, ap_enable_reg_pp0_iter135, ap_pipeline_reg_pp0_iter134_exitcond_reg_472, gmem_RVALID)
    begin
                ap_condition_1658 <= ((ap_const_lv1_1 = ap_CS_fsm_pp0_stage0) and (ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and not(((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))));
    end process;


    ap_condition_1670_assign_proc : process(ap_CS_fsm_pp1_stage0, ap_enable_reg_pp1_iter1, isIter_reg_494, ap_enable_reg_pp1_iter135, ap_pipeline_reg_pp1_iter134_exitcond9_reg_485, gmem_RVALID)
    begin
                ap_condition_1670 <= ((ap_const_lv1_1 = ap_CS_fsm_pp1_stage0) and (ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and not(((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))));
    end process;


    ap_done_assign_proc : process(ap_CS_fsm_state416, gmem_BVALID)
    begin
        if (((ap_const_lv1_1 = ap_CS_fsm_state416) and not((gmem_BVALID = ap_const_logic_0)))) then 
            ap_done <= ap_const_logic_1;
        else 
            ap_done <= ap_const_logic_0;
        end if; 
    end process;


    ap_idle_assign_proc : process(ap_start, ap_CS_fsm_state1)
    begin
        if (((ap_const_logic_0 = ap_start) and (ap_CS_fsm_state1 = ap_const_lv1_1))) then 
            ap_idle <= ap_const_logic_1;
        else 
            ap_idle <= ap_const_logic_0;
        end if; 
    end process;


    ap_ready_assign_proc : process(ap_CS_fsm_state416, gmem_BVALID)
    begin
        if (((ap_const_lv1_1 = ap_CS_fsm_state416) and not((gmem_BVALID = ap_const_logic_0)))) then 
            ap_ready <= ap_const_logic_1;
        else 
            ap_ready <= ap_const_logic_0;
        end if; 
    end process;


    ap_rst_n_inv_assign_proc : process(ap_rst_n)
    begin
                ap_rst_n_inv <= not(ap_rst_n);
    end process;


    ap_sig_ioackin_gmem_ARREADY_assign_proc : process(gmem_ARREADY, ap_reg_ioackin_gmem_ARREADY)
    begin
        if ((ap_const_logic_0 = ap_reg_ioackin_gmem_ARREADY)) then 
            ap_sig_ioackin_gmem_ARREADY <= gmem_ARREADY;
        else 
            ap_sig_ioackin_gmem_ARREADY <= ap_const_logic_1;
        end if; 
    end process;


    ap_sig_ioackin_gmem_AWREADY_assign_proc : process(gmem_AWREADY, ap_reg_ioackin_gmem_AWREADY)
    begin
        if ((ap_const_logic_0 = ap_reg_ioackin_gmem_AWREADY)) then 
            ap_sig_ioackin_gmem_AWREADY <= gmem_AWREADY;
        else 
            ap_sig_ioackin_gmem_AWREADY <= ap_const_logic_1;
        end if; 
    end process;


    ap_sig_ioackin_gmem_WREADY_assign_proc : process(gmem_WREADY, ap_reg_ioackin_gmem_WREADY)
    begin
        if ((ap_const_logic_0 = ap_reg_ioackin_gmem_WREADY)) then 
            ap_sig_ioackin_gmem_WREADY <= gmem_WREADY;
        else 
            ap_sig_ioackin_gmem_WREADY <= ap_const_logic_1;
        end if; 
    end process;

    exitcond9_fu_336_p2 <= "1" when (indvar7_phi_fu_207_p4 = ap_const_lv5_10) else "0";
    exitcond_fu_308_p2 <= "1" when (indvar_phi_fu_195_p4 = ap_const_lv5_10) else "0";

    gmem_ARADDR_assign_proc : process(arg_x_reg_455, arg_y_reg_461, ap_reg_ioackin_gmem_ARREADY, ap_condition_1658, ap_condition_1670)
    begin
        if ((ap_const_logic_0 = ap_reg_ioackin_gmem_ARREADY)) then
            if ((ap_condition_1670 = ap_const_boolean_1)) then 
                gmem_ARADDR <= arg_y_reg_461;
            elsif ((ap_condition_1658 = ap_const_boolean_1)) then 
                gmem_ARADDR <= arg_x_reg_455;
            else 
                gmem_ARADDR <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
            end if;
        else 
            gmem_ARADDR <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
        end if; 
    end process;


    gmem_ARVALID_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_enable_reg_pp0_iter1, isIter0_reg_481, ap_enable_reg_pp0_iter135, ap_pipeline_reg_pp0_iter134_exitcond_reg_472, ap_CS_fsm_pp1_stage0, ap_enable_reg_pp1_iter1, isIter_reg_494, ap_enable_reg_pp1_iter135, ap_pipeline_reg_pp1_iter134_exitcond9_reg_485, gmem_RVALID, ap_reg_ioackin_gmem_ARREADY)
    begin
        if ((((ap_const_lv1_1 = ap_CS_fsm_pp0_stage0) and (ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and not(((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))) and (ap_const_logic_0 = ap_reg_ioackin_gmem_ARREADY)) or ((ap_const_lv1_1 = ap_CS_fsm_pp1_stage0) and (ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_reg_ioackin_gmem_ARREADY) and not(((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))))) then 
            gmem_ARVALID <= ap_const_logic_1;
        else 
            gmem_ARVALID <= ap_const_logic_0;
        end if; 
    end process;


    gmem_AWVALID_assign_proc : process(ap_CS_fsm_state278, ap_reg_ioackin_gmem_AWREADY)
    begin
        if (((ap_const_lv1_1 = ap_CS_fsm_state278) and (ap_const_logic_0 = ap_reg_ioackin_gmem_AWREADY))) then 
            gmem_AWVALID <= ap_const_logic_1;
        else 
            gmem_AWVALID <= ap_const_logic_0;
        end if; 
    end process;


    gmem_BREADY_assign_proc : process(ap_CS_fsm_state416, gmem_BVALID)
    begin
        if (((ap_const_lv1_1 = ap_CS_fsm_state416) and not((gmem_BVALID = ap_const_logic_0)))) then 
            gmem_BREADY <= ap_const_logic_1;
        else 
            gmem_BREADY <= ap_const_logic_0;
        end if; 
    end process;


    gmem_RREADY_assign_proc : process(ap_enable_reg_pp0_iter1, isIter0_reg_481, ap_enable_reg_pp0_iter135, ap_pipeline_reg_pp0_iter134_exitcond_reg_472, ap_enable_reg_pp1_iter1, isIter_reg_494, ap_enable_reg_pp1_iter135, ap_pipeline_reg_pp1_iter134_exitcond9_reg_485, gmem_RVALID, ap_sig_ioackin_gmem_ARREADY)
    begin
        if ((((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0))))) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0))))))) then 
            gmem_RREADY <= ap_const_logic_1;
        else 
            gmem_RREADY <= ap_const_logic_0;
        end if; 
    end process;

    gmem_WDATA <= tmp_3_reg_536;

    gmem_WVALID_assign_proc : process(ap_CS_fsm_state285, ap_reg_ioackin_gmem_WREADY)
    begin
        if (((ap_const_lv1_1 = ap_CS_fsm_state285) and (ap_const_logic_0 = ap_reg_ioackin_gmem_WREADY))) then 
            gmem_WVALID <= ap_const_logic_1;
        else 
            gmem_WVALID <= ap_const_logic_0;
        end if; 
    end process;


    gmem_blk_n_AR_assign_proc : process(m_axi_gmem_ARREADY, ap_CS_fsm_pp0_stage0, ap_enable_reg_pp0_iter1, isIter0_reg_481, ap_CS_fsm_pp1_stage0, ap_enable_reg_pp1_iter1, isIter_reg_494)
    begin
        if ((((ap_const_lv1_1 = ap_CS_fsm_pp0_stage0) and (ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0))) or ((ap_const_lv1_1 = ap_CS_fsm_pp1_stage0) and (ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494))))) then 
            gmem_blk_n_AR <= m_axi_gmem_ARREADY;
        else 
            gmem_blk_n_AR <= ap_const_logic_1;
        end if; 
    end process;


    gmem_blk_n_AW_assign_proc : process(m_axi_gmem_AWREADY, ap_CS_fsm_state278)
    begin
        if (((ap_const_lv1_1 = ap_CS_fsm_state278))) then 
            gmem_blk_n_AW <= m_axi_gmem_AWREADY;
        else 
            gmem_blk_n_AW <= ap_const_logic_1;
        end if; 
    end process;


    gmem_blk_n_B_assign_proc : process(m_axi_gmem_BVALID, ap_CS_fsm_state416)
    begin
        if (((ap_const_lv1_1 = ap_CS_fsm_state416))) then 
            gmem_blk_n_B <= m_axi_gmem_BVALID;
        else 
            gmem_blk_n_B <= ap_const_logic_1;
        end if; 
    end process;


    gmem_blk_n_R_assign_proc : process(m_axi_gmem_RVALID, ap_enable_reg_pp0_iter135, ap_pipeline_reg_pp0_iter134_exitcond_reg_472, ap_enable_reg_pp1_iter135, ap_pipeline_reg_pp1_iter134_exitcond9_reg_485)
    begin
        if ((((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485)))) then 
            gmem_blk_n_R <= m_axi_gmem_RVALID;
        else 
            gmem_blk_n_R <= ap_const_logic_1;
        end if; 
    end process;


    gmem_blk_n_W_assign_proc : process(m_axi_gmem_WREADY, ap_CS_fsm_state285)
    begin
        if (((ap_const_lv1_1 = ap_CS_fsm_state285))) then 
            gmem_blk_n_W <= m_axi_gmem_WREADY;
        else 
            gmem_blk_n_W <= ap_const_logic_1;
        end if; 
    end process;

    indvar7_cast_fu_354_p1 <= std_logic_vector(resize(unsigned(ap_pipeline_reg_pp1_iter135_indvar7_reg_203),32));

    indvar7_phi_fu_207_p4_assign_proc : process(ap_CS_fsm_pp1_stage0, ap_enable_reg_pp1_iter1, exitcond9_reg_485, indvar7_reg_203, indvar_next8_reg_489)
    begin
        if (((ap_const_lv1_1 = ap_CS_fsm_pp1_stage0) and (ap_const_logic_1 = ap_enable_reg_pp1_iter1) and (ap_const_lv1_0 = exitcond9_reg_485))) then 
            indvar7_phi_fu_207_p4 <= indvar_next8_reg_489;
        else 
            indvar7_phi_fu_207_p4 <= indvar7_reg_203;
        end if; 
    end process;

    indvar_cast_fu_326_p1 <= std_logic_vector(resize(unsigned(ap_pipeline_reg_pp0_iter135_indvar_reg_191),32));
    indvar_inc_reg2mem_fu_405_p2 <= std_logic_vector(unsigned(indvar_reg2mem44_0_i_reg_215) + unsigned(ap_const_lv5_1));
    indvar_next8_fu_342_p2 <= std_logic_vector(unsigned(indvar7_phi_fu_207_p4) + unsigned(ap_const_lv5_1));
    indvar_next_fu_314_p2 <= std_logic_vector(unsigned(indvar_phi_fu_195_p4) + unsigned(ap_const_lv5_1));

    indvar_phi_fu_195_p4_assign_proc : process(ap_CS_fsm_pp0_stage0, ap_enable_reg_pp0_iter1, exitcond_reg_472, indvar_reg_191, indvar_next_reg_476)
    begin
        if (((ap_const_lv1_1 = ap_CS_fsm_pp0_stage0) and (ap_const_logic_1 = ap_enable_reg_pp0_iter1) and (ap_const_lv1_0 = exitcond_reg_472))) then 
            indvar_phi_fu_195_p4 <= indvar_next_reg_476;
        else 
            indvar_phi_fu_195_p4 <= indvar_reg_191;
        end if; 
    end process;

    indvar_reg2mem44_0_i_1_fu_411_p1 <= std_logic_vector(resize(unsigned(indvar_reg2mem44_0_i_reg_215),6));
    isIter0_fu_320_p2 <= "1" when (indvar_phi_fu_195_p4 = ap_const_lv5_0) else "0";
    isIter_fu_348_p2 <= "1" when (indvar7_phi_fu_207_p4 = ap_const_lv5_0) else "0";
    tmp1_fu_415_p2 <= std_logic_vector(unsigned(indvar_reg2mem44_0_i_1_fu_411_p1) + unsigned(tmp_cast_reg_450));
    tmp_10_fu_264_p1 <= std_logic_vector(resize(unsigned(tmp_4_fu_254_p4),32));
    tmp_11_fu_284_p1 <= std_logic_vector(resize(unsigned(tmp_5_fu_274_p4),32));
    tmp_12_fu_294_p4 <= z(31 downto 2);
    tmp_13_fu_371_p1 <= global_offset_x_read_reg_435(30 - 1 downto 0);
    tmp_14_fu_374_p2 <= std_logic_vector(unsigned(tmp_7_fu_364_p3) + unsigned(tmp_13_fu_371_p1));
    tmp_15_fu_380_p1 <= std_logic_vector(resize(unsigned(tmp_14_fu_374_p2),31));
    tmp_16_fu_384_p2 <= std_logic_vector(unsigned(tmp_6_cast_reg_467) + unsigned(tmp_15_fu_380_p1));
    tmp_17_fu_389_p1 <= std_logic_vector(resize(unsigned(tmp_16_reg_498),32));
    tmp_1_fu_238_p1 <= group_id_x(26 - 1 downto 0);
    tmp_2_cast1_fu_425_p1 <= std_logic_vector(resize(unsigned(tmp_2_fu_420_p2),32));
    tmp_2_fu_420_p2 <= std_logic_vector(unsigned(tmp_reg_440) + unsigned(tmp1_fu_415_p2));
    tmp_4_fu_254_p4 <= x(31 downto 2);
    tmp_5_fu_274_p4 <= y(31 downto 2);
    tmp_6_cast_fu_304_p1 <= std_logic_vector(resize(unsigned(tmp_12_fu_294_p4),31));
    tmp_6_fu_242_p1 <= group_id_x(2 - 1 downto 0);
    tmp_7_fu_364_p3 <= (tmp_1_reg_445 & ap_const_lv4_0);
    tmp_9_fu_399_p2 <= "1" when (indvar_reg2mem44_0_i_reg_215 = ap_const_lv5_10) else "0";
    tmp_cast_fu_246_p3 <= (tmp_6_fu_242_p1 & ap_const_lv4_0);
    tmp_fu_234_p1 <= global_offset_x(6 - 1 downto 0);

    x0_address0_assign_proc : process(ap_CS_fsm_state279, ap_enable_reg_pp0_iter136, indvar_cast_fu_326_p1, tmp_2_cast1_fu_425_p1)
    begin
        if (((ap_const_lv1_1 = ap_CS_fsm_state279))) then 
            x0_address0 <= tmp_2_cast1_fu_425_p1(4 - 1 downto 0);
        elsif ((ap_const_logic_1 = ap_enable_reg_pp0_iter136)) then 
            x0_address0 <= indvar_cast_fu_326_p1(4 - 1 downto 0);
        else 
            x0_address0 <= "XXXX";
        end if; 
    end process;


    x0_ce0_assign_proc : process(ap_enable_reg_pp0_iter1, isIter0_reg_481, ap_enable_reg_pp0_iter135, ap_pipeline_reg_pp0_iter134_exitcond_reg_472, gmem_RVALID, ap_sig_ioackin_gmem_ARREADY, ap_CS_fsm_state279, ap_enable_reg_pp0_iter136)
    begin
        if ((((ap_const_lv1_1 = ap_CS_fsm_state279)) or (not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp0_iter136)))) then 
            x0_ce0 <= ap_const_logic_1;
        else 
            x0_ce0 <= ap_const_logic_0;
        end if; 
    end process;

    x0_d0 <= reg_230;

    x0_we0_assign_proc : process(ap_enable_reg_pp0_iter1, isIter0_reg_481, ap_enable_reg_pp0_iter135, ap_pipeline_reg_pp0_iter134_exitcond_reg_472, gmem_RVALID, ap_sig_ioackin_gmem_ARREADY, ap_pipeline_reg_pp0_iter135_exitcond_reg_472, ap_enable_reg_pp0_iter136)
    begin
        if (((not((((ap_const_logic_1 = ap_enable_reg_pp0_iter1) and not((isIter0_reg_481 = ap_const_lv1_0)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp0_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter134_exitcond_reg_472) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp0_iter136) and (ap_const_lv1_0 = ap_pipeline_reg_pp0_iter135_exitcond_reg_472)))) then 
            x0_we0 <= ap_const_logic_1;
        else 
            x0_we0 <= ap_const_logic_0;
        end if; 
    end process;


    y0_address0_assign_proc : process(ap_CS_fsm_state279, ap_enable_reg_pp1_iter136, indvar7_cast_fu_354_p1, tmp_2_cast1_fu_425_p1)
    begin
        if (((ap_const_lv1_1 = ap_CS_fsm_state279))) then 
            y0_address0 <= tmp_2_cast1_fu_425_p1(4 - 1 downto 0);
        elsif ((ap_const_logic_1 = ap_enable_reg_pp1_iter136)) then 
            y0_address0 <= indvar7_cast_fu_354_p1(4 - 1 downto 0);
        else 
            y0_address0 <= "XXXX";
        end if; 
    end process;


    y0_ce0_assign_proc : process(ap_enable_reg_pp1_iter1, isIter_reg_494, ap_enable_reg_pp1_iter135, ap_pipeline_reg_pp1_iter134_exitcond9_reg_485, gmem_RVALID, ap_sig_ioackin_gmem_ARREADY, ap_CS_fsm_state279, ap_enable_reg_pp1_iter136)
    begin
        if ((((ap_const_lv1_1 = ap_CS_fsm_state279)) or (not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp1_iter136)))) then 
            y0_ce0 <= ap_const_logic_1;
        else 
            y0_ce0 <= ap_const_logic_0;
        end if; 
    end process;

    y0_d0 <= reg_230;

    y0_we0_assign_proc : process(ap_enable_reg_pp1_iter1, isIter_reg_494, ap_enable_reg_pp1_iter135, ap_pipeline_reg_pp1_iter134_exitcond9_reg_485, gmem_RVALID, ap_sig_ioackin_gmem_ARREADY, ap_pipeline_reg_pp1_iter135_exitcond9_reg_485, ap_enable_reg_pp1_iter136)
    begin
        if (((not((((ap_const_logic_1 = ap_enable_reg_pp1_iter1) and not((ap_const_lv1_0 = isIter_reg_494)) and (ap_const_logic_0 = ap_sig_ioackin_gmem_ARREADY)) or ((ap_const_logic_1 = ap_enable_reg_pp1_iter135) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter134_exitcond9_reg_485) and (gmem_RVALID = ap_const_logic_0)))) and (ap_const_logic_1 = ap_enable_reg_pp1_iter136) and (ap_const_lv1_0 = ap_pipeline_reg_pp1_iter135_exitcond9_reg_485)))) then 
            y0_we0 <= ap_const_logic_1;
        else 
            y0_we0 <= ap_const_logic_0;
        end if; 
    end process;

end behav;
